
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom1 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom1 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2d",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"2a"),
    10 => (x"fd",x"00",x"4f",x"4f"),
    11 => (x"d4",x"ee",x"c2",x"87"),
    12 => (x"86",x"c0",x"c6",x"4e"),
    13 => (x"49",x"d4",x"ee",x"c2"),
    14 => (x"48",x"f4",x"db",x"c2"),
    15 => (x"40",x"40",x"c0",x"89"),
    16 => (x"89",x"d0",x"40",x"40"),
    17 => (x"c1",x"87",x"f6",x"03"),
    18 => (x"00",x"87",x"df",x"db"),
    19 => (x"1e",x"87",x"fc",x"98"),
    20 => (x"1e",x"73",x"1e",x"72"),
    21 => (x"02",x"11",x"48",x"12"),
    22 => (x"c3",x"4b",x"87",x"ca"),
    23 => (x"73",x"9b",x"98",x"df"),
    24 => (x"87",x"f0",x"02",x"88"),
    25 => (x"4a",x"26",x"4b",x"26"),
    26 => (x"73",x"1e",x"4f",x"26"),
    27 => (x"c1",x"1e",x"72",x"1e"),
    28 => (x"87",x"ca",x"04",x"8b"),
    29 => (x"02",x"11",x"48",x"12"),
    30 => (x"02",x"88",x"87",x"c4"),
    31 => (x"4a",x"26",x"87",x"f1"),
    32 => (x"4f",x"26",x"4b",x"26"),
    33 => (x"73",x"1e",x"74",x"1e"),
    34 => (x"c1",x"1e",x"72",x"1e"),
    35 => (x"87",x"d0",x"04",x"8b"),
    36 => (x"02",x"11",x"48",x"12"),
    37 => (x"c3",x"4c",x"87",x"ca"),
    38 => (x"74",x"9c",x"98",x"df"),
    39 => (x"87",x"eb",x"02",x"88"),
    40 => (x"4b",x"26",x"4a",x"26"),
    41 => (x"4f",x"26",x"4c",x"26"),
    42 => (x"81",x"48",x"73",x"1e"),
    43 => (x"c5",x"02",x"a9",x"73"),
    44 => (x"05",x"53",x"12",x"87"),
    45 => (x"4f",x"26",x"87",x"f6"),
    46 => (x"4a",x"66",x"c4",x"1e"),
    47 => (x"51",x"12",x"48",x"71"),
    48 => (x"26",x"87",x"fb",x"05"),
    49 => (x"66",x"c4",x"1e",x"4f"),
    50 => (x"ff",x"48",x"11",x"4a"),
    51 => (x"c1",x"78",x"08",x"d4"),
    52 => (x"87",x"f5",x"05",x"8a"),
    53 => (x"c4",x"1e",x"4f",x"26"),
    54 => (x"d4",x"ff",x"4a",x"66"),
    55 => (x"78",x"ff",x"c3",x"48"),
    56 => (x"8a",x"c1",x"51",x"68"),
    57 => (x"26",x"87",x"f3",x"05"),
    58 => (x"1e",x"73",x"1e",x"4f"),
    59 => (x"c3",x"4b",x"d4",x"ff"),
    60 => (x"4a",x"6b",x"7b",x"ff"),
    61 => (x"6b",x"7b",x"ff",x"c3"),
    62 => (x"72",x"32",x"c8",x"49"),
    63 => (x"7b",x"ff",x"c3",x"b1"),
    64 => (x"31",x"c8",x"4a",x"6b"),
    65 => (x"ff",x"c3",x"b2",x"71"),
    66 => (x"c8",x"49",x"6b",x"7b"),
    67 => (x"71",x"b1",x"72",x"32"),
    68 => (x"26",x"87",x"c4",x"48"),
    69 => (x"26",x"4c",x"26",x"4d"),
    70 => (x"0e",x"4f",x"26",x"4b"),
    71 => (x"5d",x"5c",x"5b",x"5e"),
    72 => (x"ff",x"4a",x"71",x"0e"),
    73 => (x"49",x"72",x"4c",x"d4"),
    74 => (x"71",x"99",x"ff",x"c3"),
    75 => (x"f4",x"db",x"c2",x"7c"),
    76 => (x"87",x"c8",x"05",x"bf"),
    77 => (x"c9",x"48",x"66",x"d0"),
    78 => (x"58",x"a6",x"d4",x"30"),
    79 => (x"d8",x"49",x"66",x"d0"),
    80 => (x"99",x"ff",x"c3",x"29"),
    81 => (x"66",x"d0",x"7c",x"71"),
    82 => (x"c3",x"29",x"d0",x"49"),
    83 => (x"7c",x"71",x"99",x"ff"),
    84 => (x"c8",x"49",x"66",x"d0"),
    85 => (x"99",x"ff",x"c3",x"29"),
    86 => (x"66",x"d0",x"7c",x"71"),
    87 => (x"99",x"ff",x"c3",x"49"),
    88 => (x"49",x"72",x"7c",x"71"),
    89 => (x"ff",x"c3",x"29",x"d0"),
    90 => (x"6c",x"7c",x"71",x"99"),
    91 => (x"ff",x"f0",x"c9",x"4b"),
    92 => (x"ab",x"ff",x"c3",x"4d"),
    93 => (x"c3",x"87",x"d0",x"05"),
    94 => (x"4b",x"6c",x"7c",x"ff"),
    95 => (x"c6",x"02",x"8d",x"c1"),
    96 => (x"ab",x"ff",x"c3",x"87"),
    97 => (x"73",x"87",x"f0",x"02"),
    98 => (x"87",x"c7",x"fe",x"48"),
    99 => (x"ff",x"49",x"c0",x"1e"),
   100 => (x"ff",x"c3",x"48",x"d4"),
   101 => (x"c3",x"81",x"c1",x"78"),
   102 => (x"04",x"a9",x"b7",x"c8"),
   103 => (x"4f",x"26",x"87",x"f1"),
   104 => (x"e7",x"1e",x"73",x"1e"),
   105 => (x"df",x"f8",x"c4",x"87"),
   106 => (x"c0",x"1e",x"c0",x"4b"),
   107 => (x"f7",x"c1",x"f0",x"ff"),
   108 => (x"87",x"e7",x"fd",x"49"),
   109 => (x"a8",x"c1",x"86",x"c4"),
   110 => (x"87",x"ea",x"c0",x"05"),
   111 => (x"c3",x"48",x"d4",x"ff"),
   112 => (x"c0",x"c1",x"78",x"ff"),
   113 => (x"c0",x"c0",x"c0",x"c0"),
   114 => (x"f0",x"e1",x"c0",x"1e"),
   115 => (x"fd",x"49",x"e9",x"c1"),
   116 => (x"86",x"c4",x"87",x"c9"),
   117 => (x"ca",x"05",x"98",x"70"),
   118 => (x"48",x"d4",x"ff",x"87"),
   119 => (x"c1",x"78",x"ff",x"c3"),
   120 => (x"fe",x"87",x"cb",x"48"),
   121 => (x"8b",x"c1",x"87",x"e6"),
   122 => (x"87",x"fd",x"fe",x"05"),
   123 => (x"e6",x"fc",x"48",x"c0"),
   124 => (x"1e",x"73",x"1e",x"87"),
   125 => (x"c3",x"48",x"d4",x"ff"),
   126 => (x"4b",x"d3",x"78",x"ff"),
   127 => (x"ff",x"c0",x"1e",x"c0"),
   128 => (x"49",x"c1",x"c1",x"f0"),
   129 => (x"c4",x"87",x"d4",x"fc"),
   130 => (x"05",x"98",x"70",x"86"),
   131 => (x"d4",x"ff",x"87",x"ca"),
   132 => (x"78",x"ff",x"c3",x"48"),
   133 => (x"87",x"cb",x"48",x"c1"),
   134 => (x"c1",x"87",x"f1",x"fd"),
   135 => (x"db",x"ff",x"05",x"8b"),
   136 => (x"fb",x"48",x"c0",x"87"),
   137 => (x"5e",x"0e",x"87",x"f1"),
   138 => (x"ff",x"0e",x"5c",x"5b"),
   139 => (x"db",x"fd",x"4c",x"d4"),
   140 => (x"1e",x"ea",x"c6",x"87"),
   141 => (x"c1",x"f0",x"e1",x"c0"),
   142 => (x"de",x"fb",x"49",x"c8"),
   143 => (x"c1",x"86",x"c4",x"87"),
   144 => (x"87",x"c8",x"02",x"a8"),
   145 => (x"c0",x"87",x"ea",x"fe"),
   146 => (x"87",x"e2",x"c1",x"48"),
   147 => (x"70",x"87",x"da",x"fa"),
   148 => (x"ff",x"ff",x"cf",x"49"),
   149 => (x"a9",x"ea",x"c6",x"99"),
   150 => (x"fe",x"87",x"c8",x"02"),
   151 => (x"48",x"c0",x"87",x"d3"),
   152 => (x"c3",x"87",x"cb",x"c1"),
   153 => (x"f1",x"c0",x"7c",x"ff"),
   154 => (x"87",x"f4",x"fc",x"4b"),
   155 => (x"c0",x"02",x"98",x"70"),
   156 => (x"1e",x"c0",x"87",x"eb"),
   157 => (x"c1",x"f0",x"ff",x"c0"),
   158 => (x"de",x"fa",x"49",x"fa"),
   159 => (x"70",x"86",x"c4",x"87"),
   160 => (x"87",x"d9",x"05",x"98"),
   161 => (x"6c",x"7c",x"ff",x"c3"),
   162 => (x"7c",x"ff",x"c3",x"49"),
   163 => (x"c1",x"7c",x"7c",x"7c"),
   164 => (x"c4",x"02",x"99",x"c0"),
   165 => (x"d5",x"48",x"c1",x"87"),
   166 => (x"d1",x"48",x"c0",x"87"),
   167 => (x"05",x"ab",x"c2",x"87"),
   168 => (x"48",x"c0",x"87",x"c4"),
   169 => (x"8b",x"c1",x"87",x"c8"),
   170 => (x"87",x"fd",x"fe",x"05"),
   171 => (x"e4",x"f9",x"48",x"c0"),
   172 => (x"1e",x"73",x"1e",x"87"),
   173 => (x"48",x"f4",x"db",x"c2"),
   174 => (x"4b",x"c7",x"78",x"c1"),
   175 => (x"c2",x"48",x"d0",x"ff"),
   176 => (x"87",x"c8",x"fb",x"78"),
   177 => (x"c3",x"48",x"d0",x"ff"),
   178 => (x"c0",x"1e",x"c0",x"78"),
   179 => (x"c0",x"c1",x"d0",x"e5"),
   180 => (x"87",x"c7",x"f9",x"49"),
   181 => (x"a8",x"c1",x"86",x"c4"),
   182 => (x"4b",x"87",x"c1",x"05"),
   183 => (x"c5",x"05",x"ab",x"c2"),
   184 => (x"c0",x"48",x"c0",x"87"),
   185 => (x"8b",x"c1",x"87",x"f9"),
   186 => (x"87",x"d0",x"ff",x"05"),
   187 => (x"c2",x"87",x"f7",x"fc"),
   188 => (x"70",x"58",x"f8",x"db"),
   189 => (x"87",x"cd",x"05",x"98"),
   190 => (x"ff",x"c0",x"1e",x"c1"),
   191 => (x"49",x"d0",x"c1",x"f0"),
   192 => (x"c4",x"87",x"d8",x"f8"),
   193 => (x"48",x"d4",x"ff",x"86"),
   194 => (x"c4",x"78",x"ff",x"c3"),
   195 => (x"db",x"c2",x"87",x"e0"),
   196 => (x"d0",x"ff",x"58",x"fc"),
   197 => (x"ff",x"78",x"c2",x"48"),
   198 => (x"ff",x"c3",x"48",x"d4"),
   199 => (x"f7",x"48",x"c1",x"78"),
   200 => (x"5e",x"0e",x"87",x"f5"),
   201 => (x"0e",x"5d",x"5c",x"5b"),
   202 => (x"ff",x"c3",x"4a",x"71"),
   203 => (x"4c",x"d4",x"ff",x"4d"),
   204 => (x"d0",x"ff",x"7c",x"75"),
   205 => (x"78",x"c3",x"c4",x"48"),
   206 => (x"1e",x"72",x"7c",x"75"),
   207 => (x"c1",x"f0",x"ff",x"c0"),
   208 => (x"d6",x"f7",x"49",x"d8"),
   209 => (x"70",x"86",x"c4",x"87"),
   210 => (x"87",x"c5",x"02",x"98"),
   211 => (x"f0",x"c0",x"48",x"c0"),
   212 => (x"c3",x"7c",x"75",x"87"),
   213 => (x"c0",x"c8",x"7c",x"fe"),
   214 => (x"49",x"66",x"d4",x"1e"),
   215 => (x"c4",x"87",x"e6",x"f5"),
   216 => (x"75",x"7c",x"75",x"86"),
   217 => (x"d8",x"7c",x"75",x"7c"),
   218 => (x"75",x"4b",x"e0",x"da"),
   219 => (x"99",x"49",x"6c",x"7c"),
   220 => (x"c1",x"87",x"c5",x"05"),
   221 => (x"87",x"f3",x"05",x"8b"),
   222 => (x"d0",x"ff",x"7c",x"75"),
   223 => (x"c1",x"78",x"c2",x"48"),
   224 => (x"87",x"cf",x"f6",x"48"),
   225 => (x"4a",x"d4",x"ff",x"1e"),
   226 => (x"c4",x"48",x"d0",x"ff"),
   227 => (x"ff",x"c3",x"78",x"d1"),
   228 => (x"05",x"89",x"c1",x"7a"),
   229 => (x"4f",x"26",x"87",x"f8"),
   230 => (x"71",x"1e",x"73",x"1e"),
   231 => (x"cd",x"ee",x"c5",x"4b"),
   232 => (x"d4",x"ff",x"4a",x"df"),
   233 => (x"78",x"ff",x"c3",x"48"),
   234 => (x"fe",x"c3",x"48",x"68"),
   235 => (x"87",x"c5",x"02",x"a8"),
   236 => (x"ed",x"05",x"8a",x"c1"),
   237 => (x"05",x"9a",x"72",x"87"),
   238 => (x"48",x"c0",x"87",x"c5"),
   239 => (x"73",x"87",x"ea",x"c0"),
   240 => (x"87",x"cc",x"02",x"9b"),
   241 => (x"73",x"1e",x"66",x"c8"),
   242 => (x"87",x"ca",x"f4",x"49"),
   243 => (x"87",x"c6",x"86",x"c4"),
   244 => (x"fe",x"49",x"66",x"c8"),
   245 => (x"d4",x"ff",x"87",x"ee"),
   246 => (x"78",x"ff",x"c3",x"48"),
   247 => (x"05",x"9b",x"73",x"78"),
   248 => (x"d0",x"ff",x"87",x"c5"),
   249 => (x"c1",x"78",x"d0",x"48"),
   250 => (x"87",x"eb",x"f4",x"48"),
   251 => (x"71",x"1e",x"73",x"1e"),
   252 => (x"ff",x"4b",x"c0",x"4a"),
   253 => (x"ff",x"c3",x"48",x"d4"),
   254 => (x"48",x"d0",x"ff",x"78"),
   255 => (x"ff",x"78",x"c3",x"c4"),
   256 => (x"ff",x"c3",x"48",x"d4"),
   257 => (x"c0",x"1e",x"72",x"78"),
   258 => (x"d1",x"c1",x"f0",x"ff"),
   259 => (x"87",x"cb",x"f4",x"49"),
   260 => (x"98",x"70",x"86",x"c4"),
   261 => (x"c8",x"87",x"cd",x"05"),
   262 => (x"66",x"cc",x"1e",x"c0"),
   263 => (x"87",x"f8",x"fd",x"49"),
   264 => (x"4b",x"70",x"86",x"c4"),
   265 => (x"c2",x"48",x"d0",x"ff"),
   266 => (x"f3",x"48",x"73",x"78"),
   267 => (x"5e",x"0e",x"87",x"e9"),
   268 => (x"0e",x"5d",x"5c",x"5b"),
   269 => (x"ff",x"c0",x"1e",x"c0"),
   270 => (x"49",x"c9",x"c1",x"f0"),
   271 => (x"d2",x"87",x"dc",x"f3"),
   272 => (x"fc",x"db",x"c2",x"1e"),
   273 => (x"87",x"d0",x"fd",x"49"),
   274 => (x"4c",x"c0",x"86",x"c8"),
   275 => (x"b7",x"d2",x"84",x"c1"),
   276 => (x"87",x"f8",x"04",x"ac"),
   277 => (x"97",x"fc",x"db",x"c2"),
   278 => (x"c0",x"c3",x"49",x"bf"),
   279 => (x"a9",x"c0",x"c1",x"99"),
   280 => (x"87",x"e7",x"c0",x"05"),
   281 => (x"97",x"c3",x"dc",x"c2"),
   282 => (x"31",x"d0",x"49",x"bf"),
   283 => (x"97",x"c4",x"dc",x"c2"),
   284 => (x"32",x"c8",x"4a",x"bf"),
   285 => (x"dc",x"c2",x"b1",x"72"),
   286 => (x"4a",x"bf",x"97",x"c5"),
   287 => (x"cf",x"4c",x"71",x"b1"),
   288 => (x"9c",x"ff",x"ff",x"ff"),
   289 => (x"34",x"ca",x"84",x"c1"),
   290 => (x"c2",x"87",x"e7",x"c1"),
   291 => (x"bf",x"97",x"c5",x"dc"),
   292 => (x"c6",x"31",x"c1",x"49"),
   293 => (x"c6",x"dc",x"c2",x"99"),
   294 => (x"c7",x"4a",x"bf",x"97"),
   295 => (x"b1",x"72",x"2a",x"b7"),
   296 => (x"97",x"c1",x"dc",x"c2"),
   297 => (x"cf",x"4d",x"4a",x"bf"),
   298 => (x"c2",x"dc",x"c2",x"9d"),
   299 => (x"c3",x"4a",x"bf",x"97"),
   300 => (x"c2",x"32",x"ca",x"9a"),
   301 => (x"bf",x"97",x"c3",x"dc"),
   302 => (x"73",x"33",x"c2",x"4b"),
   303 => (x"c4",x"dc",x"c2",x"b2"),
   304 => (x"c3",x"4b",x"bf",x"97"),
   305 => (x"b7",x"c6",x"9b",x"c0"),
   306 => (x"c2",x"b2",x"73",x"2b"),
   307 => (x"71",x"48",x"c1",x"81"),
   308 => (x"c1",x"49",x"70",x"30"),
   309 => (x"70",x"30",x"75",x"48"),
   310 => (x"c1",x"4c",x"72",x"4d"),
   311 => (x"c8",x"94",x"71",x"84"),
   312 => (x"06",x"ad",x"b7",x"c0"),
   313 => (x"34",x"c1",x"87",x"cc"),
   314 => (x"c0",x"c8",x"2d",x"b7"),
   315 => (x"ff",x"01",x"ad",x"b7"),
   316 => (x"48",x"74",x"87",x"f4"),
   317 => (x"0e",x"87",x"dc",x"f0"),
   318 => (x"5d",x"5c",x"5b",x"5e"),
   319 => (x"c2",x"86",x"f8",x"0e"),
   320 => (x"c0",x"48",x"e2",x"e4"),
   321 => (x"da",x"dc",x"c2",x"78"),
   322 => (x"fb",x"49",x"c0",x"1e"),
   323 => (x"86",x"c4",x"87",x"de"),
   324 => (x"c5",x"05",x"98",x"70"),
   325 => (x"c9",x"48",x"c0",x"87"),
   326 => (x"4d",x"c0",x"87",x"ce"),
   327 => (x"f2",x"c0",x"7e",x"c1"),
   328 => (x"c2",x"49",x"bf",x"c1"),
   329 => (x"71",x"4a",x"d0",x"dd"),
   330 => (x"fd",x"ec",x"4b",x"c8"),
   331 => (x"05",x"98",x"70",x"87"),
   332 => (x"7e",x"c0",x"87",x"c2"),
   333 => (x"bf",x"fd",x"f1",x"c0"),
   334 => (x"ec",x"dd",x"c2",x"49"),
   335 => (x"4b",x"c8",x"71",x"4a"),
   336 => (x"70",x"87",x"e7",x"ec"),
   337 => (x"87",x"c2",x"05",x"98"),
   338 => (x"02",x"6e",x"7e",x"c0"),
   339 => (x"c2",x"87",x"fd",x"c0"),
   340 => (x"4d",x"bf",x"e0",x"e3"),
   341 => (x"9f",x"d8",x"e4",x"c2"),
   342 => (x"c5",x"48",x"7e",x"bf"),
   343 => (x"05",x"a8",x"ea",x"d6"),
   344 => (x"e3",x"c2",x"87",x"c7"),
   345 => (x"ce",x"4d",x"bf",x"e0"),
   346 => (x"ca",x"48",x"6e",x"87"),
   347 => (x"02",x"a8",x"d5",x"e9"),
   348 => (x"48",x"c0",x"87",x"c5"),
   349 => (x"c2",x"87",x"f1",x"c7"),
   350 => (x"75",x"1e",x"da",x"dc"),
   351 => (x"87",x"ec",x"f9",x"49"),
   352 => (x"98",x"70",x"86",x"c4"),
   353 => (x"c0",x"87",x"c5",x"05"),
   354 => (x"87",x"dc",x"c7",x"48"),
   355 => (x"bf",x"fd",x"f1",x"c0"),
   356 => (x"ec",x"dd",x"c2",x"49"),
   357 => (x"4b",x"c8",x"71",x"4a"),
   358 => (x"70",x"87",x"cf",x"eb"),
   359 => (x"87",x"c8",x"05",x"98"),
   360 => (x"48",x"e2",x"e4",x"c2"),
   361 => (x"87",x"da",x"78",x"c1"),
   362 => (x"bf",x"c1",x"f2",x"c0"),
   363 => (x"d0",x"dd",x"c2",x"49"),
   364 => (x"4b",x"c8",x"71",x"4a"),
   365 => (x"70",x"87",x"f3",x"ea"),
   366 => (x"c5",x"c0",x"02",x"98"),
   367 => (x"c6",x"48",x"c0",x"87"),
   368 => (x"e4",x"c2",x"87",x"e6"),
   369 => (x"49",x"bf",x"97",x"d8"),
   370 => (x"05",x"a9",x"d5",x"c1"),
   371 => (x"c2",x"87",x"cd",x"c0"),
   372 => (x"bf",x"97",x"d9",x"e4"),
   373 => (x"a9",x"ea",x"c2",x"49"),
   374 => (x"87",x"c5",x"c0",x"02"),
   375 => (x"c7",x"c6",x"48",x"c0"),
   376 => (x"da",x"dc",x"c2",x"87"),
   377 => (x"48",x"7e",x"bf",x"97"),
   378 => (x"02",x"a8",x"e9",x"c3"),
   379 => (x"6e",x"87",x"ce",x"c0"),
   380 => (x"a8",x"eb",x"c3",x"48"),
   381 => (x"87",x"c5",x"c0",x"02"),
   382 => (x"eb",x"c5",x"48",x"c0"),
   383 => (x"e5",x"dc",x"c2",x"87"),
   384 => (x"99",x"49",x"bf",x"97"),
   385 => (x"87",x"cc",x"c0",x"05"),
   386 => (x"97",x"e6",x"dc",x"c2"),
   387 => (x"a9",x"c2",x"49",x"bf"),
   388 => (x"87",x"c5",x"c0",x"02"),
   389 => (x"cf",x"c5",x"48",x"c0"),
   390 => (x"e7",x"dc",x"c2",x"87"),
   391 => (x"c2",x"48",x"bf",x"97"),
   392 => (x"70",x"58",x"de",x"e4"),
   393 => (x"88",x"c1",x"48",x"4c"),
   394 => (x"58",x"e2",x"e4",x"c2"),
   395 => (x"97",x"e8",x"dc",x"c2"),
   396 => (x"81",x"75",x"49",x"bf"),
   397 => (x"97",x"e9",x"dc",x"c2"),
   398 => (x"32",x"c8",x"4a",x"bf"),
   399 => (x"c2",x"7e",x"a1",x"72"),
   400 => (x"6e",x"48",x"ef",x"e8"),
   401 => (x"ea",x"dc",x"c2",x"78"),
   402 => (x"c8",x"48",x"bf",x"97"),
   403 => (x"e4",x"c2",x"58",x"a6"),
   404 => (x"c2",x"02",x"bf",x"e2"),
   405 => (x"f1",x"c0",x"87",x"d4"),
   406 => (x"c2",x"49",x"bf",x"fd"),
   407 => (x"71",x"4a",x"ec",x"dd"),
   408 => (x"c5",x"e8",x"4b",x"c8"),
   409 => (x"02",x"98",x"70",x"87"),
   410 => (x"c0",x"87",x"c5",x"c0"),
   411 => (x"87",x"f8",x"c3",x"48"),
   412 => (x"bf",x"da",x"e4",x"c2"),
   413 => (x"c3",x"e9",x"c2",x"4c"),
   414 => (x"ff",x"dc",x"c2",x"5c"),
   415 => (x"c8",x"49",x"bf",x"97"),
   416 => (x"fe",x"dc",x"c2",x"31"),
   417 => (x"a1",x"4a",x"bf",x"97"),
   418 => (x"c0",x"dd",x"c2",x"49"),
   419 => (x"d0",x"4a",x"bf",x"97"),
   420 => (x"49",x"a1",x"72",x"32"),
   421 => (x"97",x"c1",x"dd",x"c2"),
   422 => (x"32",x"d8",x"4a",x"bf"),
   423 => (x"c4",x"49",x"a1",x"72"),
   424 => (x"e8",x"c2",x"91",x"66"),
   425 => (x"c2",x"81",x"bf",x"ef"),
   426 => (x"c2",x"59",x"f7",x"e8"),
   427 => (x"bf",x"97",x"c7",x"dd"),
   428 => (x"c2",x"32",x"c8",x"4a"),
   429 => (x"bf",x"97",x"c6",x"dd"),
   430 => (x"c2",x"4a",x"a2",x"4b"),
   431 => (x"bf",x"97",x"c8",x"dd"),
   432 => (x"73",x"33",x"d0",x"4b"),
   433 => (x"dd",x"c2",x"4a",x"a2"),
   434 => (x"4b",x"bf",x"97",x"c9"),
   435 => (x"33",x"d8",x"9b",x"cf"),
   436 => (x"c2",x"4a",x"a2",x"73"),
   437 => (x"c2",x"5a",x"fb",x"e8"),
   438 => (x"4a",x"bf",x"f7",x"e8"),
   439 => (x"92",x"74",x"8a",x"c2"),
   440 => (x"48",x"fb",x"e8",x"c2"),
   441 => (x"c1",x"78",x"a1",x"72"),
   442 => (x"dc",x"c2",x"87",x"ca"),
   443 => (x"49",x"bf",x"97",x"ec"),
   444 => (x"dc",x"c2",x"31",x"c8"),
   445 => (x"4a",x"bf",x"97",x"eb"),
   446 => (x"e4",x"c2",x"49",x"a1"),
   447 => (x"e4",x"c2",x"59",x"ea"),
   448 => (x"c5",x"49",x"bf",x"e6"),
   449 => (x"81",x"ff",x"c7",x"31"),
   450 => (x"e9",x"c2",x"29",x"c9"),
   451 => (x"dc",x"c2",x"59",x"c3"),
   452 => (x"4a",x"bf",x"97",x"f1"),
   453 => (x"dc",x"c2",x"32",x"c8"),
   454 => (x"4b",x"bf",x"97",x"f0"),
   455 => (x"66",x"c4",x"4a",x"a2"),
   456 => (x"c2",x"82",x"6e",x"92"),
   457 => (x"c2",x"5a",x"ff",x"e8"),
   458 => (x"c0",x"48",x"f7",x"e8"),
   459 => (x"f3",x"e8",x"c2",x"78"),
   460 => (x"78",x"a1",x"72",x"48"),
   461 => (x"48",x"c3",x"e9",x"c2"),
   462 => (x"bf",x"f7",x"e8",x"c2"),
   463 => (x"c7",x"e9",x"c2",x"78"),
   464 => (x"fb",x"e8",x"c2",x"48"),
   465 => (x"e4",x"c2",x"78",x"bf"),
   466 => (x"c0",x"02",x"bf",x"e2"),
   467 => (x"48",x"74",x"87",x"c9"),
   468 => (x"7e",x"70",x"30",x"c4"),
   469 => (x"c2",x"87",x"c9",x"c0"),
   470 => (x"48",x"bf",x"ff",x"e8"),
   471 => (x"7e",x"70",x"30",x"c4"),
   472 => (x"48",x"e6",x"e4",x"c2"),
   473 => (x"48",x"c1",x"78",x"6e"),
   474 => (x"4d",x"26",x"8e",x"f8"),
   475 => (x"4b",x"26",x"4c",x"26"),
   476 => (x"5e",x"0e",x"4f",x"26"),
   477 => (x"0e",x"5d",x"5c",x"5b"),
   478 => (x"e4",x"c2",x"4a",x"71"),
   479 => (x"cb",x"02",x"bf",x"e2"),
   480 => (x"c7",x"4b",x"72",x"87"),
   481 => (x"c1",x"4c",x"72",x"2b"),
   482 => (x"87",x"c9",x"9c",x"ff"),
   483 => (x"2b",x"c8",x"4b",x"72"),
   484 => (x"ff",x"c3",x"4c",x"72"),
   485 => (x"ef",x"e8",x"c2",x"9c"),
   486 => (x"f1",x"c0",x"83",x"bf"),
   487 => (x"02",x"ab",x"bf",x"f9"),
   488 => (x"f1",x"c0",x"87",x"d9"),
   489 => (x"dc",x"c2",x"5b",x"fd"),
   490 => (x"49",x"73",x"1e",x"da"),
   491 => (x"c4",x"87",x"fd",x"f0"),
   492 => (x"05",x"98",x"70",x"86"),
   493 => (x"48",x"c0",x"87",x"c5"),
   494 => (x"c2",x"87",x"e6",x"c0"),
   495 => (x"02",x"bf",x"e2",x"e4"),
   496 => (x"49",x"74",x"87",x"d2"),
   497 => (x"dc",x"c2",x"91",x"c4"),
   498 => (x"4d",x"69",x"81",x"da"),
   499 => (x"ff",x"ff",x"ff",x"cf"),
   500 => (x"87",x"cb",x"9d",x"ff"),
   501 => (x"91",x"c2",x"49",x"74"),
   502 => (x"81",x"da",x"dc",x"c2"),
   503 => (x"75",x"4d",x"69",x"9f"),
   504 => (x"87",x"c6",x"fe",x"48"),
   505 => (x"5c",x"5b",x"5e",x"0e"),
   506 => (x"71",x"1e",x"0e",x"5d"),
   507 => (x"c1",x"1e",x"c0",x"4d"),
   508 => (x"87",x"ee",x"ca",x"49"),
   509 => (x"4c",x"70",x"86",x"c4"),
   510 => (x"c0",x"c1",x"02",x"9c"),
   511 => (x"ea",x"e4",x"c2",x"87"),
   512 => (x"e1",x"49",x"75",x"4a"),
   513 => (x"98",x"70",x"87",x"c9"),
   514 => (x"87",x"f1",x"c0",x"02"),
   515 => (x"49",x"75",x"4a",x"74"),
   516 => (x"ef",x"e1",x"4b",x"cb"),
   517 => (x"02",x"98",x"70",x"87"),
   518 => (x"c0",x"87",x"e2",x"c0"),
   519 => (x"02",x"9c",x"74",x"1e"),
   520 => (x"a6",x"c4",x"87",x"c7"),
   521 => (x"c5",x"78",x"c0",x"48"),
   522 => (x"48",x"a6",x"c4",x"87"),
   523 => (x"66",x"c4",x"78",x"c1"),
   524 => (x"87",x"ee",x"c9",x"49"),
   525 => (x"4c",x"70",x"86",x"c4"),
   526 => (x"c0",x"ff",x"05",x"9c"),
   527 => (x"26",x"48",x"74",x"87"),
   528 => (x"0e",x"87",x"e7",x"fc"),
   529 => (x"5d",x"5c",x"5b",x"5e"),
   530 => (x"4b",x"71",x"1e",x"0e"),
   531 => (x"87",x"c5",x"05",x"9b"),
   532 => (x"e5",x"c1",x"48",x"c0"),
   533 => (x"4d",x"a3",x"c8",x"87"),
   534 => (x"66",x"d4",x"7d",x"c0"),
   535 => (x"d4",x"87",x"c7",x"02"),
   536 => (x"05",x"bf",x"97",x"66"),
   537 => (x"48",x"c0",x"87",x"c5"),
   538 => (x"d4",x"87",x"cf",x"c1"),
   539 => (x"f3",x"fd",x"49",x"66"),
   540 => (x"9c",x"4c",x"70",x"87"),
   541 => (x"87",x"c0",x"c1",x"02"),
   542 => (x"69",x"49",x"a4",x"dc"),
   543 => (x"49",x"a4",x"da",x"7d"),
   544 => (x"9f",x"4a",x"a3",x"c4"),
   545 => (x"e4",x"c2",x"7a",x"69"),
   546 => (x"d2",x"02",x"bf",x"e2"),
   547 => (x"49",x"a4",x"d4",x"87"),
   548 => (x"c0",x"49",x"69",x"9f"),
   549 => (x"71",x"99",x"ff",x"ff"),
   550 => (x"70",x"30",x"d0",x"48"),
   551 => (x"c0",x"87",x"c2",x"7e"),
   552 => (x"48",x"49",x"6e",x"7e"),
   553 => (x"7a",x"70",x"80",x"6a"),
   554 => (x"a3",x"cc",x"7b",x"c0"),
   555 => (x"d0",x"79",x"6a",x"49"),
   556 => (x"79",x"c0",x"49",x"a3"),
   557 => (x"87",x"c2",x"48",x"74"),
   558 => (x"fa",x"26",x"48",x"c0"),
   559 => (x"5e",x"0e",x"87",x"ec"),
   560 => (x"0e",x"5d",x"5c",x"5b"),
   561 => (x"f1",x"c0",x"4c",x"71"),
   562 => (x"78",x"ff",x"48",x"f9"),
   563 => (x"c1",x"02",x"9c",x"74"),
   564 => (x"a4",x"c8",x"87",x"ca"),
   565 => (x"c1",x"02",x"69",x"49"),
   566 => (x"66",x"d0",x"87",x"c2"),
   567 => (x"82",x"49",x"6c",x"4a"),
   568 => (x"d0",x"5a",x"a6",x"d4"),
   569 => (x"c2",x"b9",x"4d",x"66"),
   570 => (x"4a",x"bf",x"de",x"e4"),
   571 => (x"99",x"72",x"ba",x"ff"),
   572 => (x"c0",x"02",x"99",x"71"),
   573 => (x"a4",x"c4",x"87",x"e4"),
   574 => (x"f9",x"49",x"6b",x"4b"),
   575 => (x"7b",x"70",x"87",x"f4"),
   576 => (x"bf",x"da",x"e4",x"c2"),
   577 => (x"71",x"81",x"6c",x"49"),
   578 => (x"c2",x"b9",x"75",x"7c"),
   579 => (x"4a",x"bf",x"de",x"e4"),
   580 => (x"99",x"72",x"ba",x"ff"),
   581 => (x"ff",x"05",x"99",x"71"),
   582 => (x"7c",x"75",x"87",x"dc"),
   583 => (x"1e",x"87",x"cb",x"f9"),
   584 => (x"4b",x"71",x"1e",x"73"),
   585 => (x"87",x"c7",x"02",x"9b"),
   586 => (x"69",x"49",x"a3",x"c8"),
   587 => (x"c0",x"87",x"c5",x"05"),
   588 => (x"87",x"eb",x"c0",x"48"),
   589 => (x"bf",x"f3",x"e8",x"c2"),
   590 => (x"49",x"a3",x"c4",x"4a"),
   591 => (x"89",x"c2",x"49",x"69"),
   592 => (x"bf",x"da",x"e4",x"c2"),
   593 => (x"4a",x"a2",x"71",x"91"),
   594 => (x"bf",x"de",x"e4",x"c2"),
   595 => (x"71",x"99",x"6b",x"49"),
   596 => (x"66",x"c8",x"4a",x"a2"),
   597 => (x"ea",x"49",x"72",x"1e"),
   598 => (x"86",x"c4",x"87",x"d2"),
   599 => (x"f8",x"48",x"49",x"70"),
   600 => (x"73",x"1e",x"87",x"cc"),
   601 => (x"9b",x"4b",x"71",x"1e"),
   602 => (x"c8",x"87",x"c7",x"02"),
   603 => (x"05",x"69",x"49",x"a3"),
   604 => (x"48",x"c0",x"87",x"c5"),
   605 => (x"c2",x"87",x"eb",x"c0"),
   606 => (x"4a",x"bf",x"f3",x"e8"),
   607 => (x"69",x"49",x"a3",x"c4"),
   608 => (x"c2",x"89",x"c2",x"49"),
   609 => (x"91",x"bf",x"da",x"e4"),
   610 => (x"c2",x"4a",x"a2",x"71"),
   611 => (x"49",x"bf",x"de",x"e4"),
   612 => (x"a2",x"71",x"99",x"6b"),
   613 => (x"1e",x"66",x"c8",x"4a"),
   614 => (x"c5",x"e6",x"49",x"72"),
   615 => (x"70",x"86",x"c4",x"87"),
   616 => (x"c9",x"f7",x"48",x"49"),
   617 => (x"5b",x"5e",x"0e",x"87"),
   618 => (x"1e",x"0e",x"5d",x"5c"),
   619 => (x"66",x"d4",x"4b",x"71"),
   620 => (x"73",x"2c",x"c9",x"4c"),
   621 => (x"cf",x"c1",x"02",x"9b"),
   622 => (x"49",x"a3",x"c8",x"87"),
   623 => (x"c7",x"c1",x"02",x"69"),
   624 => (x"4d",x"a3",x"d0",x"87"),
   625 => (x"c2",x"7d",x"66",x"d4"),
   626 => (x"49",x"bf",x"de",x"e4"),
   627 => (x"4a",x"6b",x"b9",x"ff"),
   628 => (x"ac",x"71",x"7e",x"99"),
   629 => (x"c0",x"87",x"cd",x"03"),
   630 => (x"a3",x"cc",x"7d",x"7b"),
   631 => (x"49",x"a3",x"c4",x"4a"),
   632 => (x"87",x"c2",x"79",x"6a"),
   633 => (x"9c",x"74",x"8c",x"72"),
   634 => (x"49",x"87",x"dd",x"02"),
   635 => (x"fb",x"49",x"73",x"1e"),
   636 => (x"86",x"c4",x"87",x"cc"),
   637 => (x"c7",x"49",x"66",x"d4"),
   638 => (x"cb",x"02",x"99",x"ff"),
   639 => (x"da",x"dc",x"c2",x"87"),
   640 => (x"fc",x"49",x"73",x"1e"),
   641 => (x"86",x"c4",x"87",x"d9"),
   642 => (x"87",x"de",x"f5",x"26"),
   643 => (x"71",x"1e",x"73",x"1e"),
   644 => (x"c0",x"02",x"9b",x"4b"),
   645 => (x"e9",x"c2",x"87",x"e4"),
   646 => (x"4a",x"73",x"5b",x"c7"),
   647 => (x"e4",x"c2",x"8a",x"c2"),
   648 => (x"92",x"49",x"bf",x"da"),
   649 => (x"bf",x"f3",x"e8",x"c2"),
   650 => (x"c2",x"80",x"72",x"48"),
   651 => (x"71",x"58",x"cb",x"e9"),
   652 => (x"c2",x"30",x"c4",x"48"),
   653 => (x"c0",x"58",x"ea",x"e4"),
   654 => (x"e9",x"c2",x"87",x"ed"),
   655 => (x"e8",x"c2",x"48",x"c3"),
   656 => (x"c2",x"78",x"bf",x"f7"),
   657 => (x"c2",x"48",x"c7",x"e9"),
   658 => (x"78",x"bf",x"fb",x"e8"),
   659 => (x"bf",x"e2",x"e4",x"c2"),
   660 => (x"c2",x"87",x"c9",x"02"),
   661 => (x"49",x"bf",x"da",x"e4"),
   662 => (x"87",x"c7",x"31",x"c4"),
   663 => (x"bf",x"ff",x"e8",x"c2"),
   664 => (x"c2",x"31",x"c4",x"49"),
   665 => (x"f4",x"59",x"ea",x"e4"),
   666 => (x"5e",x"0e",x"87",x"c4"),
   667 => (x"71",x"0e",x"5c",x"5b"),
   668 => (x"72",x"4b",x"c0",x"4a"),
   669 => (x"e1",x"c0",x"02",x"9a"),
   670 => (x"49",x"a2",x"da",x"87"),
   671 => (x"c2",x"4b",x"69",x"9f"),
   672 => (x"02",x"bf",x"e2",x"e4"),
   673 => (x"a2",x"d4",x"87",x"cf"),
   674 => (x"49",x"69",x"9f",x"49"),
   675 => (x"ff",x"ff",x"c0",x"4c"),
   676 => (x"c2",x"34",x"d0",x"9c"),
   677 => (x"74",x"4c",x"c0",x"87"),
   678 => (x"49",x"73",x"b3",x"49"),
   679 => (x"f3",x"87",x"ed",x"fd"),
   680 => (x"5e",x"0e",x"87",x"ca"),
   681 => (x"0e",x"5d",x"5c",x"5b"),
   682 => (x"4a",x"71",x"86",x"f4"),
   683 => (x"9a",x"72",x"7e",x"c0"),
   684 => (x"c2",x"87",x"d8",x"02"),
   685 => (x"c0",x"48",x"d6",x"dc"),
   686 => (x"ce",x"dc",x"c2",x"78"),
   687 => (x"c7",x"e9",x"c2",x"48"),
   688 => (x"dc",x"c2",x"78",x"bf"),
   689 => (x"e9",x"c2",x"48",x"d2"),
   690 => (x"c2",x"78",x"bf",x"c3"),
   691 => (x"c0",x"48",x"f7",x"e4"),
   692 => (x"e6",x"e4",x"c2",x"50"),
   693 => (x"dc",x"c2",x"49",x"bf"),
   694 => (x"71",x"4a",x"bf",x"d6"),
   695 => (x"ff",x"c3",x"03",x"aa"),
   696 => (x"cf",x"49",x"72",x"87"),
   697 => (x"e0",x"c0",x"05",x"99"),
   698 => (x"da",x"dc",x"c2",x"87"),
   699 => (x"ce",x"dc",x"c2",x"1e"),
   700 => (x"dc",x"c2",x"49",x"bf"),
   701 => (x"a1",x"c1",x"48",x"ce"),
   702 => (x"ef",x"e3",x"71",x"78"),
   703 => (x"c0",x"86",x"c4",x"87"),
   704 => (x"c2",x"48",x"f5",x"f1"),
   705 => (x"cc",x"78",x"da",x"dc"),
   706 => (x"f5",x"f1",x"c0",x"87"),
   707 => (x"e0",x"c0",x"48",x"bf"),
   708 => (x"f9",x"f1",x"c0",x"80"),
   709 => (x"d6",x"dc",x"c2",x"58"),
   710 => (x"80",x"c1",x"48",x"bf"),
   711 => (x"58",x"da",x"dc",x"c2"),
   712 => (x"00",x"0c",x"75",x"27"),
   713 => (x"bf",x"97",x"bf",x"00"),
   714 => (x"c2",x"02",x"9d",x"4d"),
   715 => (x"e5",x"c3",x"87",x"e2"),
   716 => (x"db",x"c2",x"02",x"ad"),
   717 => (x"f5",x"f1",x"c0",x"87"),
   718 => (x"a3",x"cb",x"4b",x"bf"),
   719 => (x"cf",x"4c",x"11",x"49"),
   720 => (x"d2",x"c1",x"05",x"ac"),
   721 => (x"df",x"49",x"75",x"87"),
   722 => (x"cd",x"89",x"c1",x"99"),
   723 => (x"ea",x"e4",x"c2",x"91"),
   724 => (x"4a",x"a3",x"c1",x"81"),
   725 => (x"a3",x"c3",x"51",x"12"),
   726 => (x"c5",x"51",x"12",x"4a"),
   727 => (x"51",x"12",x"4a",x"a3"),
   728 => (x"12",x"4a",x"a3",x"c7"),
   729 => (x"4a",x"a3",x"c9",x"51"),
   730 => (x"a3",x"ce",x"51",x"12"),
   731 => (x"d0",x"51",x"12",x"4a"),
   732 => (x"51",x"12",x"4a",x"a3"),
   733 => (x"12",x"4a",x"a3",x"d2"),
   734 => (x"4a",x"a3",x"d4",x"51"),
   735 => (x"a3",x"d6",x"51",x"12"),
   736 => (x"d8",x"51",x"12",x"4a"),
   737 => (x"51",x"12",x"4a",x"a3"),
   738 => (x"12",x"4a",x"a3",x"dc"),
   739 => (x"4a",x"a3",x"de",x"51"),
   740 => (x"7e",x"c1",x"51",x"12"),
   741 => (x"74",x"87",x"f9",x"c0"),
   742 => (x"05",x"99",x"c8",x"49"),
   743 => (x"74",x"87",x"ea",x"c0"),
   744 => (x"05",x"99",x"d0",x"49"),
   745 => (x"66",x"dc",x"87",x"d0"),
   746 => (x"87",x"ca",x"c0",x"02"),
   747 => (x"66",x"dc",x"49",x"73"),
   748 => (x"02",x"98",x"70",x"0f"),
   749 => (x"05",x"6e",x"87",x"d3"),
   750 => (x"c2",x"87",x"c6",x"c0"),
   751 => (x"c0",x"48",x"ea",x"e4"),
   752 => (x"f5",x"f1",x"c0",x"50"),
   753 => (x"e7",x"c2",x"48",x"bf"),
   754 => (x"f7",x"e4",x"c2",x"87"),
   755 => (x"7e",x"50",x"c0",x"48"),
   756 => (x"bf",x"e6",x"e4",x"c2"),
   757 => (x"d6",x"dc",x"c2",x"49"),
   758 => (x"aa",x"71",x"4a",x"bf"),
   759 => (x"87",x"c1",x"fc",x"04"),
   760 => (x"bf",x"c7",x"e9",x"c2"),
   761 => (x"87",x"c8",x"c0",x"05"),
   762 => (x"bf",x"e2",x"e4",x"c2"),
   763 => (x"87",x"fe",x"c1",x"02"),
   764 => (x"48",x"f9",x"f1",x"c0"),
   765 => (x"dc",x"c2",x"78",x"ff"),
   766 => (x"ed",x"49",x"bf",x"d2"),
   767 => (x"49",x"70",x"87",x"f4"),
   768 => (x"59",x"d6",x"dc",x"c2"),
   769 => (x"c2",x"48",x"a6",x"c4"),
   770 => (x"78",x"bf",x"d2",x"dc"),
   771 => (x"bf",x"e2",x"e4",x"c2"),
   772 => (x"87",x"d8",x"c0",x"02"),
   773 => (x"cf",x"49",x"66",x"c4"),
   774 => (x"f8",x"ff",x"ff",x"ff"),
   775 => (x"c0",x"02",x"a9",x"99"),
   776 => (x"4d",x"c0",x"87",x"c5"),
   777 => (x"c1",x"87",x"e1",x"c0"),
   778 => (x"87",x"dc",x"c0",x"4d"),
   779 => (x"cf",x"49",x"66",x"c4"),
   780 => (x"a9",x"99",x"f8",x"ff"),
   781 => (x"87",x"c8",x"c0",x"02"),
   782 => (x"c0",x"48",x"a6",x"c8"),
   783 => (x"87",x"c5",x"c0",x"78"),
   784 => (x"c1",x"48",x"a6",x"c8"),
   785 => (x"4d",x"66",x"c8",x"78"),
   786 => (x"c0",x"05",x"9d",x"75"),
   787 => (x"66",x"c4",x"87",x"e0"),
   788 => (x"c2",x"89",x"c2",x"49"),
   789 => (x"4a",x"bf",x"da",x"e4"),
   790 => (x"f3",x"e8",x"c2",x"91"),
   791 => (x"dc",x"c2",x"4a",x"bf"),
   792 => (x"a1",x"72",x"48",x"ce"),
   793 => (x"d6",x"dc",x"c2",x"78"),
   794 => (x"f9",x"78",x"c0",x"48"),
   795 => (x"48",x"c0",x"87",x"e3"),
   796 => (x"f5",x"eb",x"8e",x"f4"),
   797 => (x"00",x"00",x"00",x"87"),
   798 => (x"ff",x"ff",x"ff",x"00"),
   799 => (x"00",x"0c",x"85",x"ff"),
   800 => (x"00",x"0c",x"8e",x"00"),
   801 => (x"54",x"41",x"46",x"00"),
   802 => (x"20",x"20",x"32",x"33"),
   803 => (x"41",x"46",x"00",x"20"),
   804 => (x"20",x"36",x"31",x"54"),
   805 => (x"1e",x"00",x"20",x"20"),
   806 => (x"c3",x"48",x"d4",x"ff"),
   807 => (x"48",x"68",x"78",x"ff"),
   808 => (x"ff",x"1e",x"4f",x"26"),
   809 => (x"ff",x"c3",x"48",x"d4"),
   810 => (x"48",x"d0",x"ff",x"78"),
   811 => (x"ff",x"78",x"e1",x"c8"),
   812 => (x"78",x"d4",x"48",x"d4"),
   813 => (x"48",x"cb",x"e9",x"c2"),
   814 => (x"50",x"bf",x"d4",x"ff"),
   815 => (x"ff",x"1e",x"4f",x"26"),
   816 => (x"e0",x"c0",x"48",x"d0"),
   817 => (x"1e",x"4f",x"26",x"78"),
   818 => (x"70",x"87",x"cc",x"ff"),
   819 => (x"c6",x"02",x"99",x"49"),
   820 => (x"a9",x"fb",x"c0",x"87"),
   821 => (x"71",x"87",x"f1",x"05"),
   822 => (x"0e",x"4f",x"26",x"48"),
   823 => (x"0e",x"5c",x"5b",x"5e"),
   824 => (x"4c",x"c0",x"4b",x"71"),
   825 => (x"70",x"87",x"f0",x"fe"),
   826 => (x"c0",x"02",x"99",x"49"),
   827 => (x"ec",x"c0",x"87",x"f9"),
   828 => (x"f2",x"c0",x"02",x"a9"),
   829 => (x"a9",x"fb",x"c0",x"87"),
   830 => (x"87",x"eb",x"c0",x"02"),
   831 => (x"ac",x"b7",x"66",x"cc"),
   832 => (x"d0",x"87",x"c7",x"03"),
   833 => (x"87",x"c2",x"02",x"66"),
   834 => (x"99",x"71",x"53",x"71"),
   835 => (x"c1",x"87",x"c2",x"02"),
   836 => (x"87",x"c3",x"fe",x"84"),
   837 => (x"02",x"99",x"49",x"70"),
   838 => (x"ec",x"c0",x"87",x"cd"),
   839 => (x"87",x"c7",x"02",x"a9"),
   840 => (x"05",x"a9",x"fb",x"c0"),
   841 => (x"d0",x"87",x"d5",x"ff"),
   842 => (x"87",x"c3",x"02",x"66"),
   843 => (x"c0",x"7b",x"97",x"c0"),
   844 => (x"c4",x"05",x"a9",x"ec"),
   845 => (x"c5",x"4a",x"74",x"87"),
   846 => (x"c0",x"4a",x"74",x"87"),
   847 => (x"48",x"72",x"8a",x"0a"),
   848 => (x"4d",x"26",x"87",x"c2"),
   849 => (x"4b",x"26",x"4c",x"26"),
   850 => (x"fd",x"1e",x"4f",x"26"),
   851 => (x"49",x"70",x"87",x"c9"),
   852 => (x"a9",x"b7",x"f0",x"c0"),
   853 => (x"c0",x"87",x"ca",x"04"),
   854 => (x"01",x"a9",x"b7",x"f9"),
   855 => (x"f0",x"c0",x"87",x"c3"),
   856 => (x"b7",x"c1",x"c1",x"89"),
   857 => (x"87",x"ca",x"04",x"a9"),
   858 => (x"a9",x"b7",x"da",x"c1"),
   859 => (x"c0",x"87",x"c3",x"01"),
   860 => (x"48",x"71",x"89",x"f7"),
   861 => (x"5e",x"0e",x"4f",x"26"),
   862 => (x"71",x"0e",x"5c",x"5b"),
   863 => (x"4c",x"d4",x"ff",x"4a"),
   864 => (x"ea",x"c0",x"49",x"72"),
   865 => (x"9b",x"4b",x"70",x"87"),
   866 => (x"c1",x"87",x"c2",x"02"),
   867 => (x"48",x"d0",x"ff",x"8b"),
   868 => (x"c1",x"78",x"c5",x"c8"),
   869 => (x"49",x"73",x"7c",x"d5"),
   870 => (x"da",x"c2",x"31",x"c6"),
   871 => (x"4a",x"bf",x"97",x"de"),
   872 => (x"70",x"b0",x"71",x"48"),
   873 => (x"48",x"d0",x"ff",x"7c"),
   874 => (x"48",x"73",x"78",x"c4"),
   875 => (x"0e",x"87",x"d5",x"fe"),
   876 => (x"5d",x"5c",x"5b",x"5e"),
   877 => (x"71",x"86",x"f8",x"0e"),
   878 => (x"fb",x"7e",x"c0",x"4c"),
   879 => (x"4b",x"c0",x"87",x"e4"),
   880 => (x"97",x"dc",x"f9",x"c0"),
   881 => (x"a9",x"c0",x"49",x"bf"),
   882 => (x"fb",x"87",x"cf",x"04"),
   883 => (x"83",x"c1",x"87",x"f9"),
   884 => (x"97",x"dc",x"f9",x"c0"),
   885 => (x"06",x"ab",x"49",x"bf"),
   886 => (x"f9",x"c0",x"87",x"f1"),
   887 => (x"02",x"bf",x"97",x"dc"),
   888 => (x"f2",x"fa",x"87",x"cf"),
   889 => (x"99",x"49",x"70",x"87"),
   890 => (x"c0",x"87",x"c6",x"02"),
   891 => (x"f1",x"05",x"a9",x"ec"),
   892 => (x"fa",x"4b",x"c0",x"87"),
   893 => (x"4d",x"70",x"87",x"e1"),
   894 => (x"c8",x"87",x"dc",x"fa"),
   895 => (x"d6",x"fa",x"58",x"a6"),
   896 => (x"c1",x"4a",x"70",x"87"),
   897 => (x"49",x"a4",x"c8",x"83"),
   898 => (x"ad",x"49",x"69",x"97"),
   899 => (x"c0",x"87",x"c7",x"02"),
   900 => (x"c0",x"05",x"ad",x"ff"),
   901 => (x"a4",x"c9",x"87",x"e7"),
   902 => (x"49",x"69",x"97",x"49"),
   903 => (x"02",x"a9",x"66",x"c4"),
   904 => (x"c0",x"48",x"87",x"c7"),
   905 => (x"d4",x"05",x"a8",x"ff"),
   906 => (x"49",x"a4",x"ca",x"87"),
   907 => (x"aa",x"49",x"69",x"97"),
   908 => (x"c0",x"87",x"c6",x"02"),
   909 => (x"c4",x"05",x"aa",x"ff"),
   910 => (x"d0",x"7e",x"c1",x"87"),
   911 => (x"ad",x"ec",x"c0",x"87"),
   912 => (x"c0",x"87",x"c6",x"02"),
   913 => (x"c4",x"05",x"ad",x"fb"),
   914 => (x"c1",x"4b",x"c0",x"87"),
   915 => (x"fe",x"02",x"6e",x"7e"),
   916 => (x"e9",x"f9",x"87",x"e1"),
   917 => (x"f8",x"48",x"73",x"87"),
   918 => (x"87",x"e6",x"fb",x"8e"),
   919 => (x"5b",x"5e",x"0e",x"00"),
   920 => (x"1e",x"0e",x"5d",x"5c"),
   921 => (x"4c",x"c0",x"4b",x"71"),
   922 => (x"c0",x"04",x"ab",x"4d"),
   923 => (x"f6",x"c0",x"87",x"e8"),
   924 => (x"9d",x"75",x"1e",x"ef"),
   925 => (x"c0",x"87",x"c4",x"02"),
   926 => (x"c1",x"87",x"c2",x"4a"),
   927 => (x"f0",x"49",x"72",x"4a"),
   928 => (x"86",x"c4",x"87",x"e0"),
   929 => (x"84",x"c1",x"7e",x"70"),
   930 => (x"87",x"c2",x"05",x"6e"),
   931 => (x"85",x"c1",x"4c",x"73"),
   932 => (x"ff",x"06",x"ac",x"73"),
   933 => (x"48",x"6e",x"87",x"d8"),
   934 => (x"26",x"4d",x"26",x"26"),
   935 => (x"26",x"4b",x"26",x"4c"),
   936 => (x"5b",x"5e",x"0e",x"4f"),
   937 => (x"1e",x"0e",x"5d",x"5c"),
   938 => (x"de",x"49",x"4c",x"71"),
   939 => (x"e5",x"e9",x"c2",x"91"),
   940 => (x"97",x"85",x"71",x"4d"),
   941 => (x"dd",x"c1",x"02",x"6d"),
   942 => (x"d0",x"e9",x"c2",x"87"),
   943 => (x"82",x"74",x"4a",x"bf"),
   944 => (x"d8",x"fe",x"49",x"72"),
   945 => (x"6e",x"7e",x"70",x"87"),
   946 => (x"87",x"f3",x"c0",x"02"),
   947 => (x"4b",x"d8",x"e9",x"c2"),
   948 => (x"49",x"cb",x"4a",x"6e"),
   949 => (x"87",x"d0",x"c7",x"ff"),
   950 => (x"93",x"cb",x"4b",x"74"),
   951 => (x"83",x"ce",x"dd",x"c1"),
   952 => (x"fc",x"c0",x"83",x"c4"),
   953 => (x"49",x"74",x"7b",x"da"),
   954 => (x"87",x"c9",x"c3",x"c1"),
   955 => (x"e9",x"c2",x"7b",x"75"),
   956 => (x"49",x"bf",x"97",x"e4"),
   957 => (x"d8",x"e9",x"c2",x"1e"),
   958 => (x"e3",x"dd",x"c1",x"49"),
   959 => (x"74",x"86",x"c4",x"87"),
   960 => (x"f0",x"c2",x"c1",x"49"),
   961 => (x"c1",x"49",x"c0",x"87"),
   962 => (x"c2",x"87",x"cf",x"c4"),
   963 => (x"c0",x"48",x"cc",x"e9"),
   964 => (x"dd",x"49",x"c1",x"78"),
   965 => (x"fd",x"26",x"87",x"cb"),
   966 => (x"6f",x"4c",x"87",x"ff"),
   967 => (x"6e",x"69",x"64",x"61"),
   968 => (x"2e",x"2e",x"2e",x"67"),
   969 => (x"5b",x"5e",x"0e",x"00"),
   970 => (x"4b",x"71",x"0e",x"5c"),
   971 => (x"d0",x"e9",x"c2",x"4a"),
   972 => (x"49",x"72",x"82",x"bf"),
   973 => (x"70",x"87",x"e6",x"fc"),
   974 => (x"c4",x"02",x"9c",x"4c"),
   975 => (x"e9",x"ec",x"49",x"87"),
   976 => (x"d0",x"e9",x"c2",x"87"),
   977 => (x"c1",x"78",x"c0",x"48"),
   978 => (x"87",x"d5",x"dc",x"49"),
   979 => (x"0e",x"87",x"cc",x"fd"),
   980 => (x"5d",x"5c",x"5b",x"5e"),
   981 => (x"c2",x"86",x"f4",x"0e"),
   982 => (x"c0",x"4d",x"da",x"dc"),
   983 => (x"48",x"a6",x"c4",x"4c"),
   984 => (x"e9",x"c2",x"78",x"c0"),
   985 => (x"c0",x"49",x"bf",x"d0"),
   986 => (x"c1",x"c1",x"06",x"a9"),
   987 => (x"da",x"dc",x"c2",x"87"),
   988 => (x"c0",x"02",x"98",x"48"),
   989 => (x"f6",x"c0",x"87",x"f8"),
   990 => (x"66",x"c8",x"1e",x"ef"),
   991 => (x"c4",x"87",x"c7",x"02"),
   992 => (x"78",x"c0",x"48",x"a6"),
   993 => (x"a6",x"c4",x"87",x"c5"),
   994 => (x"c4",x"78",x"c1",x"48"),
   995 => (x"d1",x"ec",x"49",x"66"),
   996 => (x"70",x"86",x"c4",x"87"),
   997 => (x"c4",x"84",x"c1",x"4d"),
   998 => (x"80",x"c1",x"48",x"66"),
   999 => (x"c2",x"58",x"a6",x"c8"),
  1000 => (x"49",x"bf",x"d0",x"e9"),
  1001 => (x"87",x"c6",x"03",x"ac"),
  1002 => (x"ff",x"05",x"9d",x"75"),
  1003 => (x"4c",x"c0",x"87",x"c8"),
  1004 => (x"c3",x"02",x"9d",x"75"),
  1005 => (x"f6",x"c0",x"87",x"e0"),
  1006 => (x"66",x"c8",x"1e",x"ef"),
  1007 => (x"cc",x"87",x"c7",x"02"),
  1008 => (x"78",x"c0",x"48",x"a6"),
  1009 => (x"a6",x"cc",x"87",x"c5"),
  1010 => (x"cc",x"78",x"c1",x"48"),
  1011 => (x"d1",x"eb",x"49",x"66"),
  1012 => (x"70",x"86",x"c4",x"87"),
  1013 => (x"c2",x"02",x"6e",x"7e"),
  1014 => (x"49",x"6e",x"87",x"e9"),
  1015 => (x"69",x"97",x"81",x"cb"),
  1016 => (x"02",x"99",x"d0",x"49"),
  1017 => (x"c0",x"87",x"d6",x"c1"),
  1018 => (x"74",x"4a",x"e5",x"fc"),
  1019 => (x"c1",x"91",x"cb",x"49"),
  1020 => (x"72",x"81",x"ce",x"dd"),
  1021 => (x"c3",x"81",x"c8",x"79"),
  1022 => (x"49",x"74",x"51",x"ff"),
  1023 => (x"e9",x"c2",x"91",x"de"),
  1024 => (x"85",x"71",x"4d",x"e5"),
  1025 => (x"7d",x"97",x"c1",x"c2"),
  1026 => (x"c0",x"49",x"a5",x"c1"),
  1027 => (x"e4",x"c2",x"51",x"e0"),
  1028 => (x"02",x"bf",x"97",x"ea"),
  1029 => (x"84",x"c1",x"87",x"d2"),
  1030 => (x"c2",x"4b",x"a5",x"c2"),
  1031 => (x"db",x"4a",x"ea",x"e4"),
  1032 => (x"c3",x"c2",x"ff",x"49"),
  1033 => (x"87",x"db",x"c1",x"87"),
  1034 => (x"c0",x"49",x"a5",x"cd"),
  1035 => (x"c2",x"84",x"c1",x"51"),
  1036 => (x"4a",x"6e",x"4b",x"a5"),
  1037 => (x"c1",x"ff",x"49",x"cb"),
  1038 => (x"c6",x"c1",x"87",x"ee"),
  1039 => (x"e1",x"fa",x"c0",x"87"),
  1040 => (x"cb",x"49",x"74",x"4a"),
  1041 => (x"ce",x"dd",x"c1",x"91"),
  1042 => (x"c2",x"79",x"72",x"81"),
  1043 => (x"bf",x"97",x"ea",x"e4"),
  1044 => (x"74",x"87",x"d8",x"02"),
  1045 => (x"c1",x"91",x"de",x"49"),
  1046 => (x"e5",x"e9",x"c2",x"84"),
  1047 => (x"c2",x"83",x"71",x"4b"),
  1048 => (x"dd",x"4a",x"ea",x"e4"),
  1049 => (x"ff",x"c0",x"ff",x"49"),
  1050 => (x"74",x"87",x"d8",x"87"),
  1051 => (x"c2",x"93",x"de",x"4b"),
  1052 => (x"cb",x"83",x"e5",x"e9"),
  1053 => (x"51",x"c0",x"49",x"a3"),
  1054 => (x"6e",x"73",x"84",x"c1"),
  1055 => (x"ff",x"49",x"cb",x"4a"),
  1056 => (x"c4",x"87",x"e5",x"c0"),
  1057 => (x"80",x"c1",x"48",x"66"),
  1058 => (x"c7",x"58",x"a6",x"c8"),
  1059 => (x"c5",x"c0",x"03",x"ac"),
  1060 => (x"fc",x"05",x"6e",x"87"),
  1061 => (x"48",x"74",x"87",x"e0"),
  1062 => (x"fc",x"f7",x"8e",x"f4"),
  1063 => (x"1e",x"73",x"1e",x"87"),
  1064 => (x"cb",x"49",x"4b",x"71"),
  1065 => (x"ce",x"dd",x"c1",x"91"),
  1066 => (x"4a",x"a1",x"c8",x"81"),
  1067 => (x"48",x"de",x"da",x"c2"),
  1068 => (x"a1",x"c9",x"50",x"12"),
  1069 => (x"dc",x"f9",x"c0",x"4a"),
  1070 => (x"ca",x"50",x"12",x"48"),
  1071 => (x"e4",x"e9",x"c2",x"81"),
  1072 => (x"c2",x"50",x"11",x"48"),
  1073 => (x"bf",x"97",x"e4",x"e9"),
  1074 => (x"49",x"c0",x"1e",x"49"),
  1075 => (x"87",x"d0",x"d6",x"c1"),
  1076 => (x"48",x"cc",x"e9",x"c2"),
  1077 => (x"49",x"c1",x"78",x"de"),
  1078 => (x"26",x"87",x"c6",x"d6"),
  1079 => (x"1e",x"87",x"fe",x"f6"),
  1080 => (x"cb",x"49",x"4a",x"71"),
  1081 => (x"ce",x"dd",x"c1",x"91"),
  1082 => (x"11",x"81",x"c8",x"81"),
  1083 => (x"d0",x"e9",x"c2",x"48"),
  1084 => (x"d0",x"e9",x"c2",x"58"),
  1085 => (x"c1",x"78",x"c0",x"48"),
  1086 => (x"87",x"e5",x"d5",x"49"),
  1087 => (x"c0",x"1e",x"4f",x"26"),
  1088 => (x"d5",x"fc",x"c0",x"49"),
  1089 => (x"1e",x"4f",x"26",x"87"),
  1090 => (x"d2",x"02",x"99",x"71"),
  1091 => (x"e3",x"de",x"c1",x"87"),
  1092 => (x"f7",x"50",x"c0",x"48"),
  1093 => (x"df",x"c3",x"c1",x"80"),
  1094 => (x"c7",x"dd",x"c1",x"40"),
  1095 => (x"c1",x"87",x"ce",x"78"),
  1096 => (x"c1",x"48",x"df",x"de"),
  1097 => (x"fc",x"78",x"c0",x"dd"),
  1098 => (x"fe",x"c3",x"c1",x"80"),
  1099 => (x"0e",x"4f",x"26",x"78"),
  1100 => (x"0e",x"5c",x"5b",x"5e"),
  1101 => (x"cb",x"4a",x"4c",x"71"),
  1102 => (x"ce",x"dd",x"c1",x"92"),
  1103 => (x"49",x"a2",x"c8",x"82"),
  1104 => (x"97",x"4b",x"a2",x"c9"),
  1105 => (x"97",x"1e",x"4b",x"6b"),
  1106 => (x"ca",x"1e",x"49",x"69"),
  1107 => (x"c0",x"49",x"12",x"82"),
  1108 => (x"c0",x"87",x"d0",x"e7"),
  1109 => (x"87",x"c9",x"d4",x"49"),
  1110 => (x"f9",x"c0",x"49",x"74"),
  1111 => (x"8e",x"f8",x"87",x"d7"),
  1112 => (x"1e",x"87",x"f8",x"f4"),
  1113 => (x"4b",x"71",x"1e",x"73"),
  1114 => (x"87",x"c3",x"ff",x"49"),
  1115 => (x"fe",x"fe",x"49",x"73"),
  1116 => (x"87",x"e9",x"f4",x"87"),
  1117 => (x"71",x"1e",x"73",x"1e"),
  1118 => (x"4a",x"a3",x"c6",x"4b"),
  1119 => (x"c1",x"87",x"db",x"02"),
  1120 => (x"87",x"d6",x"02",x"8a"),
  1121 => (x"da",x"c1",x"02",x"8a"),
  1122 => (x"c0",x"02",x"8a",x"87"),
  1123 => (x"02",x"8a",x"87",x"fc"),
  1124 => (x"8a",x"87",x"e1",x"c0"),
  1125 => (x"c1",x"87",x"cb",x"02"),
  1126 => (x"49",x"c7",x"87",x"db"),
  1127 => (x"c1",x"87",x"c0",x"fd"),
  1128 => (x"e9",x"c2",x"87",x"de"),
  1129 => (x"c1",x"02",x"bf",x"d0"),
  1130 => (x"c1",x"48",x"87",x"cb"),
  1131 => (x"d4",x"e9",x"c2",x"88"),
  1132 => (x"87",x"c1",x"c1",x"58"),
  1133 => (x"bf",x"d4",x"e9",x"c2"),
  1134 => (x"87",x"f9",x"c0",x"02"),
  1135 => (x"bf",x"d0",x"e9",x"c2"),
  1136 => (x"c2",x"80",x"c1",x"48"),
  1137 => (x"c0",x"58",x"d4",x"e9"),
  1138 => (x"e9",x"c2",x"87",x"eb"),
  1139 => (x"c6",x"49",x"bf",x"d0"),
  1140 => (x"d4",x"e9",x"c2",x"89"),
  1141 => (x"a9",x"b7",x"c0",x"59"),
  1142 => (x"c2",x"87",x"da",x"03"),
  1143 => (x"c0",x"48",x"d0",x"e9"),
  1144 => (x"c2",x"87",x"d2",x"78"),
  1145 => (x"02",x"bf",x"d4",x"e9"),
  1146 => (x"e9",x"c2",x"87",x"cb"),
  1147 => (x"c6",x"48",x"bf",x"d0"),
  1148 => (x"d4",x"e9",x"c2",x"80"),
  1149 => (x"d1",x"49",x"c0",x"58"),
  1150 => (x"49",x"73",x"87",x"e7"),
  1151 => (x"87",x"f5",x"f6",x"c0"),
  1152 => (x"0e",x"87",x"da",x"f2"),
  1153 => (x"0e",x"5c",x"5b",x"5e"),
  1154 => (x"66",x"cc",x"4c",x"71"),
  1155 => (x"cb",x"4b",x"74",x"1e"),
  1156 => (x"ce",x"dd",x"c1",x"93"),
  1157 => (x"4a",x"a3",x"c4",x"83"),
  1158 => (x"fa",x"fe",x"49",x"6a"),
  1159 => (x"c2",x"c1",x"87",x"da"),
  1160 => (x"a3",x"c8",x"7b",x"dd"),
  1161 => (x"51",x"66",x"d4",x"49"),
  1162 => (x"d8",x"49",x"a3",x"c9"),
  1163 => (x"a3",x"ca",x"51",x"66"),
  1164 => (x"51",x"66",x"dc",x"49"),
  1165 => (x"87",x"e3",x"f1",x"26"),
  1166 => (x"5c",x"5b",x"5e",x"0e"),
  1167 => (x"d0",x"ff",x"0e",x"5d"),
  1168 => (x"59",x"a6",x"d8",x"86"),
  1169 => (x"c0",x"48",x"a6",x"c4"),
  1170 => (x"c1",x"80",x"c4",x"78"),
  1171 => (x"c4",x"78",x"66",x"c4"),
  1172 => (x"c4",x"78",x"c1",x"80"),
  1173 => (x"c2",x"78",x"c1",x"80"),
  1174 => (x"c1",x"48",x"d4",x"e9"),
  1175 => (x"cc",x"e9",x"c2",x"78"),
  1176 => (x"a8",x"de",x"48",x"bf"),
  1177 => (x"f3",x"87",x"cb",x"05"),
  1178 => (x"49",x"70",x"87",x"e5"),
  1179 => (x"ce",x"59",x"a6",x"c8"),
  1180 => (x"ed",x"e8",x"87",x"f8"),
  1181 => (x"87",x"cf",x"e9",x"87"),
  1182 => (x"70",x"87",x"dc",x"e8"),
  1183 => (x"ac",x"fb",x"c0",x"4c"),
  1184 => (x"87",x"d0",x"c1",x"02"),
  1185 => (x"c1",x"05",x"66",x"d4"),
  1186 => (x"1e",x"c0",x"87",x"c2"),
  1187 => (x"c1",x"1e",x"c1",x"1e"),
  1188 => (x"c0",x"1e",x"c1",x"df"),
  1189 => (x"87",x"eb",x"fd",x"49"),
  1190 => (x"4a",x"66",x"d0",x"c1"),
  1191 => (x"49",x"6a",x"82",x"c4"),
  1192 => (x"51",x"74",x"81",x"c7"),
  1193 => (x"1e",x"d8",x"1e",x"c1"),
  1194 => (x"81",x"c8",x"49",x"6a"),
  1195 => (x"d8",x"87",x"ec",x"e8"),
  1196 => (x"66",x"c4",x"c1",x"86"),
  1197 => (x"01",x"a8",x"c0",x"48"),
  1198 => (x"a6",x"c4",x"87",x"c7"),
  1199 => (x"ce",x"78",x"c1",x"48"),
  1200 => (x"66",x"c4",x"c1",x"87"),
  1201 => (x"cc",x"88",x"c1",x"48"),
  1202 => (x"87",x"c3",x"58",x"a6"),
  1203 => (x"cc",x"87",x"f8",x"e7"),
  1204 => (x"78",x"c2",x"48",x"a6"),
  1205 => (x"cd",x"02",x"9c",x"74"),
  1206 => (x"66",x"c4",x"87",x"cc"),
  1207 => (x"66",x"c8",x"c1",x"48"),
  1208 => (x"c1",x"cd",x"03",x"a8"),
  1209 => (x"48",x"a6",x"d8",x"87"),
  1210 => (x"ea",x"e6",x"78",x"c0"),
  1211 => (x"c1",x"4c",x"70",x"87"),
  1212 => (x"c2",x"05",x"ac",x"d0"),
  1213 => (x"66",x"d8",x"87",x"d6"),
  1214 => (x"87",x"ce",x"e9",x"7e"),
  1215 => (x"a6",x"dc",x"49",x"70"),
  1216 => (x"87",x"d3",x"e6",x"59"),
  1217 => (x"ec",x"c0",x"4c",x"70"),
  1218 => (x"ea",x"c1",x"05",x"ac"),
  1219 => (x"49",x"66",x"c4",x"87"),
  1220 => (x"c0",x"c1",x"91",x"cb"),
  1221 => (x"a1",x"c4",x"81",x"66"),
  1222 => (x"c8",x"4d",x"6a",x"4a"),
  1223 => (x"66",x"d8",x"4a",x"a1"),
  1224 => (x"df",x"c3",x"c1",x"52"),
  1225 => (x"87",x"ef",x"e5",x"79"),
  1226 => (x"02",x"9c",x"4c",x"70"),
  1227 => (x"fb",x"c0",x"87",x"d8"),
  1228 => (x"87",x"d2",x"02",x"ac"),
  1229 => (x"de",x"e5",x"55",x"74"),
  1230 => (x"9c",x"4c",x"70",x"87"),
  1231 => (x"c0",x"87",x"c7",x"02"),
  1232 => (x"ff",x"05",x"ac",x"fb"),
  1233 => (x"e0",x"c0",x"87",x"ee"),
  1234 => (x"55",x"c1",x"c2",x"55"),
  1235 => (x"d4",x"7d",x"97",x"c0"),
  1236 => (x"a9",x"6e",x"49",x"66"),
  1237 => (x"c4",x"87",x"db",x"05"),
  1238 => (x"66",x"c8",x"48",x"66"),
  1239 => (x"87",x"ca",x"04",x"a8"),
  1240 => (x"c1",x"48",x"66",x"c4"),
  1241 => (x"58",x"a6",x"c8",x"80"),
  1242 => (x"66",x"c8",x"87",x"c8"),
  1243 => (x"cc",x"88",x"c1",x"48"),
  1244 => (x"e2",x"e4",x"58",x"a6"),
  1245 => (x"c1",x"4c",x"70",x"87"),
  1246 => (x"c8",x"05",x"ac",x"d0"),
  1247 => (x"48",x"66",x"d0",x"87"),
  1248 => (x"a6",x"d4",x"80",x"c1"),
  1249 => (x"ac",x"d0",x"c1",x"58"),
  1250 => (x"87",x"ea",x"fd",x"02"),
  1251 => (x"d4",x"48",x"a6",x"dc"),
  1252 => (x"66",x"d8",x"78",x"66"),
  1253 => (x"a8",x"66",x"dc",x"48"),
  1254 => (x"87",x"dc",x"c9",x"05"),
  1255 => (x"48",x"a6",x"e0",x"c0"),
  1256 => (x"c4",x"78",x"f0",x"c0"),
  1257 => (x"78",x"66",x"cc",x"80"),
  1258 => (x"78",x"c0",x"80",x"c4"),
  1259 => (x"c0",x"48",x"74",x"7e"),
  1260 => (x"f0",x"c0",x"88",x"fb"),
  1261 => (x"98",x"70",x"58",x"a6"),
  1262 => (x"87",x"d7",x"c8",x"02"),
  1263 => (x"c0",x"88",x"cb",x"48"),
  1264 => (x"70",x"58",x"a6",x"f0"),
  1265 => (x"e9",x"c0",x"02",x"98"),
  1266 => (x"88",x"c9",x"48",x"87"),
  1267 => (x"58",x"a6",x"f0",x"c0"),
  1268 => (x"c3",x"02",x"98",x"70"),
  1269 => (x"c4",x"48",x"87",x"e1"),
  1270 => (x"a6",x"f0",x"c0",x"88"),
  1271 => (x"02",x"98",x"70",x"58"),
  1272 => (x"c1",x"48",x"87",x"d6"),
  1273 => (x"a6",x"f0",x"c0",x"88"),
  1274 => (x"02",x"98",x"70",x"58"),
  1275 => (x"c7",x"87",x"c8",x"c3"),
  1276 => (x"e0",x"c0",x"87",x"db"),
  1277 => (x"78",x"c0",x"48",x"a6"),
  1278 => (x"c1",x"48",x"66",x"cc"),
  1279 => (x"58",x"a6",x"d0",x"80"),
  1280 => (x"70",x"87",x"d4",x"e2"),
  1281 => (x"ac",x"ec",x"c0",x"4c"),
  1282 => (x"c0",x"87",x"d5",x"02"),
  1283 => (x"c6",x"02",x"66",x"e0"),
  1284 => (x"a6",x"e4",x"c0",x"87"),
  1285 => (x"74",x"87",x"c9",x"5c"),
  1286 => (x"88",x"f0",x"c0",x"48"),
  1287 => (x"58",x"a6",x"e8",x"c0"),
  1288 => (x"02",x"ac",x"ec",x"c0"),
  1289 => (x"ee",x"e1",x"87",x"cc"),
  1290 => (x"c0",x"4c",x"70",x"87"),
  1291 => (x"ff",x"05",x"ac",x"ec"),
  1292 => (x"e0",x"c0",x"87",x"f4"),
  1293 => (x"66",x"d4",x"1e",x"66"),
  1294 => (x"ec",x"c0",x"1e",x"49"),
  1295 => (x"df",x"c1",x"1e",x"66"),
  1296 => (x"66",x"d4",x"1e",x"c1"),
  1297 => (x"87",x"fb",x"f6",x"49"),
  1298 => (x"1e",x"ca",x"1e",x"c0"),
  1299 => (x"cb",x"49",x"66",x"dc"),
  1300 => (x"66",x"d8",x"c1",x"91"),
  1301 => (x"48",x"a6",x"d8",x"81"),
  1302 => (x"d8",x"78",x"a1",x"c4"),
  1303 => (x"e1",x"49",x"bf",x"66"),
  1304 => (x"86",x"d8",x"87",x"f9"),
  1305 => (x"06",x"a8",x"b7",x"c0"),
  1306 => (x"c1",x"87",x"c7",x"c1"),
  1307 => (x"c8",x"1e",x"de",x"1e"),
  1308 => (x"e1",x"49",x"bf",x"66"),
  1309 => (x"86",x"c8",x"87",x"e5"),
  1310 => (x"c0",x"48",x"49",x"70"),
  1311 => (x"e4",x"c0",x"88",x"08"),
  1312 => (x"b7",x"c0",x"58",x"a6"),
  1313 => (x"e9",x"c0",x"06",x"a8"),
  1314 => (x"66",x"e0",x"c0",x"87"),
  1315 => (x"a8",x"b7",x"dd",x"48"),
  1316 => (x"6e",x"87",x"df",x"03"),
  1317 => (x"e0",x"c0",x"49",x"bf"),
  1318 => (x"e0",x"c0",x"81",x"66"),
  1319 => (x"c1",x"49",x"66",x"51"),
  1320 => (x"81",x"bf",x"6e",x"81"),
  1321 => (x"c0",x"51",x"c1",x"c2"),
  1322 => (x"c2",x"49",x"66",x"e0"),
  1323 => (x"81",x"bf",x"6e",x"81"),
  1324 => (x"7e",x"c1",x"51",x"c0"),
  1325 => (x"e2",x"87",x"dc",x"c4"),
  1326 => (x"e4",x"c0",x"87",x"d0"),
  1327 => (x"c9",x"e2",x"58",x"a6"),
  1328 => (x"a6",x"e8",x"c0",x"87"),
  1329 => (x"a8",x"ec",x"c0",x"58"),
  1330 => (x"87",x"cb",x"c0",x"05"),
  1331 => (x"48",x"a6",x"e4",x"c0"),
  1332 => (x"78",x"66",x"e0",x"c0"),
  1333 => (x"ff",x"87",x"c4",x"c0"),
  1334 => (x"c4",x"87",x"fc",x"de"),
  1335 => (x"91",x"cb",x"49",x"66"),
  1336 => (x"48",x"66",x"c0",x"c1"),
  1337 => (x"7e",x"70",x"80",x"71"),
  1338 => (x"82",x"c8",x"4a",x"6e"),
  1339 => (x"81",x"ca",x"49",x"6e"),
  1340 => (x"51",x"66",x"e0",x"c0"),
  1341 => (x"49",x"66",x"e4",x"c0"),
  1342 => (x"e0",x"c0",x"81",x"c1"),
  1343 => (x"48",x"c1",x"89",x"66"),
  1344 => (x"49",x"70",x"30",x"71"),
  1345 => (x"97",x"71",x"89",x"c1"),
  1346 => (x"c1",x"ed",x"c2",x"7a"),
  1347 => (x"e0",x"c0",x"49",x"bf"),
  1348 => (x"6a",x"97",x"29",x"66"),
  1349 => (x"98",x"71",x"48",x"4a"),
  1350 => (x"58",x"a6",x"f0",x"c0"),
  1351 => (x"81",x"c4",x"49",x"6e"),
  1352 => (x"66",x"dc",x"4d",x"69"),
  1353 => (x"a8",x"66",x"d8",x"48"),
  1354 => (x"87",x"c8",x"c0",x"02"),
  1355 => (x"c0",x"48",x"a6",x"d8"),
  1356 => (x"87",x"c5",x"c0",x"78"),
  1357 => (x"c1",x"48",x"a6",x"d8"),
  1358 => (x"1e",x"66",x"d8",x"78"),
  1359 => (x"75",x"1e",x"e0",x"c0"),
  1360 => (x"d6",x"de",x"ff",x"49"),
  1361 => (x"70",x"86",x"c8",x"87"),
  1362 => (x"ac",x"b7",x"c0",x"4c"),
  1363 => (x"87",x"d4",x"c1",x"06"),
  1364 => (x"e0",x"c0",x"85",x"74"),
  1365 => (x"75",x"89",x"74",x"49"),
  1366 => (x"de",x"d9",x"c1",x"4b"),
  1367 => (x"ed",x"fe",x"71",x"4a"),
  1368 => (x"85",x"c2",x"87",x"c6"),
  1369 => (x"48",x"66",x"e8",x"c0"),
  1370 => (x"ec",x"c0",x"80",x"c1"),
  1371 => (x"ec",x"c0",x"58",x"a6"),
  1372 => (x"81",x"c1",x"49",x"66"),
  1373 => (x"c0",x"02",x"a9",x"70"),
  1374 => (x"a6",x"d8",x"87",x"c8"),
  1375 => (x"c0",x"78",x"c0",x"48"),
  1376 => (x"a6",x"d8",x"87",x"c5"),
  1377 => (x"d8",x"78",x"c1",x"48"),
  1378 => (x"a4",x"c2",x"1e",x"66"),
  1379 => (x"48",x"e0",x"c0",x"49"),
  1380 => (x"49",x"70",x"88",x"71"),
  1381 => (x"ff",x"49",x"75",x"1e"),
  1382 => (x"c8",x"87",x"c0",x"dd"),
  1383 => (x"a8",x"b7",x"c0",x"86"),
  1384 => (x"87",x"c0",x"ff",x"01"),
  1385 => (x"02",x"66",x"e8",x"c0"),
  1386 => (x"6e",x"87",x"d1",x"c0"),
  1387 => (x"c0",x"81",x"c9",x"49"),
  1388 => (x"6e",x"51",x"66",x"e8"),
  1389 => (x"ef",x"c4",x"c1",x"48"),
  1390 => (x"87",x"cc",x"c0",x"78"),
  1391 => (x"81",x"c9",x"49",x"6e"),
  1392 => (x"48",x"6e",x"51",x"c2"),
  1393 => (x"78",x"e3",x"c5",x"c1"),
  1394 => (x"c6",x"c0",x"7e",x"c1"),
  1395 => (x"f6",x"db",x"ff",x"87"),
  1396 => (x"6e",x"4c",x"70",x"87"),
  1397 => (x"87",x"f5",x"c0",x"02"),
  1398 => (x"c8",x"48",x"66",x"c4"),
  1399 => (x"c0",x"04",x"a8",x"66"),
  1400 => (x"66",x"c4",x"87",x"cb"),
  1401 => (x"c8",x"80",x"c1",x"48"),
  1402 => (x"e0",x"c0",x"58",x"a6"),
  1403 => (x"48",x"66",x"c8",x"87"),
  1404 => (x"a6",x"cc",x"88",x"c1"),
  1405 => (x"87",x"d5",x"c0",x"58"),
  1406 => (x"05",x"ac",x"c6",x"c1"),
  1407 => (x"cc",x"87",x"c8",x"c0"),
  1408 => (x"80",x"c1",x"48",x"66"),
  1409 => (x"ff",x"58",x"a6",x"d0"),
  1410 => (x"70",x"87",x"fc",x"da"),
  1411 => (x"48",x"66",x"d0",x"4c"),
  1412 => (x"a6",x"d4",x"80",x"c1"),
  1413 => (x"02",x"9c",x"74",x"58"),
  1414 => (x"c4",x"87",x"cb",x"c0"),
  1415 => (x"c8",x"c1",x"48",x"66"),
  1416 => (x"f2",x"04",x"a8",x"66"),
  1417 => (x"da",x"ff",x"87",x"ff"),
  1418 => (x"66",x"c4",x"87",x"d4"),
  1419 => (x"03",x"a8",x"c7",x"48"),
  1420 => (x"c2",x"87",x"e5",x"c0"),
  1421 => (x"c0",x"48",x"d4",x"e9"),
  1422 => (x"49",x"66",x"c4",x"78"),
  1423 => (x"c0",x"c1",x"91",x"cb"),
  1424 => (x"a1",x"c4",x"81",x"66"),
  1425 => (x"c0",x"4a",x"6a",x"4a"),
  1426 => (x"66",x"c4",x"79",x"52"),
  1427 => (x"c8",x"80",x"c1",x"48"),
  1428 => (x"a8",x"c7",x"58",x"a6"),
  1429 => (x"87",x"db",x"ff",x"04"),
  1430 => (x"e0",x"8e",x"d0",x"ff"),
  1431 => (x"20",x"3a",x"87",x"fb"),
  1432 => (x"1e",x"73",x"1e",x"00"),
  1433 => (x"02",x"9b",x"4b",x"71"),
  1434 => (x"e9",x"c2",x"87",x"c6"),
  1435 => (x"78",x"c0",x"48",x"d0"),
  1436 => (x"e9",x"c2",x"1e",x"c7"),
  1437 => (x"1e",x"49",x"bf",x"d0"),
  1438 => (x"1e",x"ce",x"dd",x"c1"),
  1439 => (x"bf",x"cc",x"e9",x"c2"),
  1440 => (x"87",x"f4",x"ee",x"49"),
  1441 => (x"e9",x"c2",x"86",x"cc"),
  1442 => (x"e9",x"49",x"bf",x"cc"),
  1443 => (x"9b",x"73",x"87",x"f9"),
  1444 => (x"c1",x"87",x"c8",x"02"),
  1445 => (x"c0",x"49",x"ce",x"dd"),
  1446 => (x"ff",x"87",x"ec",x"e5"),
  1447 => (x"1e",x"87",x"fe",x"df"),
  1448 => (x"48",x"de",x"da",x"c2"),
  1449 => (x"de",x"c1",x"50",x"c0"),
  1450 => (x"c0",x"49",x"bf",x"f1"),
  1451 => (x"c0",x"87",x"c4",x"fb"),
  1452 => (x"1e",x"4f",x"26",x"48"),
  1453 => (x"c1",x"87",x"e9",x"c7"),
  1454 => (x"87",x"e5",x"fe",x"49"),
  1455 => (x"87",x"f1",x"ef",x"fe"),
  1456 => (x"cd",x"02",x"98",x"70"),
  1457 => (x"ee",x"f8",x"fe",x"87"),
  1458 => (x"02",x"98",x"70",x"87"),
  1459 => (x"4a",x"c1",x"87",x"c4"),
  1460 => (x"4a",x"c0",x"87",x"c2"),
  1461 => (x"ce",x"05",x"9a",x"72"),
  1462 => (x"c1",x"1e",x"c0",x"87"),
  1463 => (x"c0",x"49",x"c7",x"dc"),
  1464 => (x"c4",x"87",x"f3",x"f0"),
  1465 => (x"c0",x"87",x"fe",x"86"),
  1466 => (x"c0",x"87",x"dd",x"ff"),
  1467 => (x"d2",x"dc",x"c1",x"1e"),
  1468 => (x"e1",x"f0",x"c0",x"49"),
  1469 => (x"fe",x"1e",x"c0",x"87"),
  1470 => (x"49",x"70",x"87",x"e5"),
  1471 => (x"87",x"d6",x"f0",x"c0"),
  1472 => (x"f8",x"87",x"dc",x"c3"),
  1473 => (x"53",x"4f",x"26",x"8e"),
  1474 => (x"61",x"66",x"20",x"44"),
  1475 => (x"64",x"65",x"6c",x"69"),
  1476 => (x"6f",x"42",x"00",x"2e"),
  1477 => (x"6e",x"69",x"74",x"6f"),
  1478 => (x"2e",x"2e",x"2e",x"67"),
  1479 => (x"e8",x"c0",x"1e",x"00"),
  1480 => (x"f3",x"c0",x"87",x"c1"),
  1481 => (x"87",x"f6",x"87",x"e6"),
  1482 => (x"c2",x"1e",x"4f",x"26"),
  1483 => (x"c0",x"48",x"d0",x"e9"),
  1484 => (x"cc",x"e9",x"c2",x"78"),
  1485 => (x"fd",x"78",x"c0",x"48"),
  1486 => (x"87",x"e1",x"87",x"f9"),
  1487 => (x"4f",x"26",x"48",x"c0"),
  1488 => (x"78",x"45",x"20",x"80"),
  1489 => (x"80",x"00",x"74",x"69"),
  1490 => (x"63",x"61",x"42",x"20"),
  1491 => (x"10",x"df",x"00",x"6b"),
  1492 => (x"2a",x"65",x"00",x"00"),
  1493 => (x"00",x"00",x"00",x"00"),
  1494 => (x"00",x"10",x"df",x"00"),
  1495 => (x"00",x"2a",x"83",x"00"),
  1496 => (x"00",x"00",x"00",x"00"),
  1497 => (x"00",x"00",x"10",x"df"),
  1498 => (x"00",x"00",x"2a",x"a1"),
  1499 => (x"df",x"00",x"00",x"00"),
  1500 => (x"bf",x"00",x"00",x"10"),
  1501 => (x"00",x"00",x"00",x"2a"),
  1502 => (x"10",x"df",x"00",x"00"),
  1503 => (x"2a",x"dd",x"00",x"00"),
  1504 => (x"00",x"00",x"00",x"00"),
  1505 => (x"00",x"10",x"df",x"00"),
  1506 => (x"00",x"2a",x"fb",x"00"),
  1507 => (x"00",x"00",x"00",x"00"),
  1508 => (x"00",x"00",x"10",x"df"),
  1509 => (x"00",x"00",x"2b",x"19"),
  1510 => (x"df",x"00",x"00",x"00"),
  1511 => (x"00",x"00",x"00",x"10"),
  1512 => (x"00",x"00",x"00",x"00"),
  1513 => (x"11",x"74",x"00",x"00"),
  1514 => (x"00",x"00",x"00",x"00"),
  1515 => (x"00",x"00",x"00",x"00"),
  1516 => (x"00",x"17",x"b5",x"00"),
  1517 => (x"4f",x"4f",x"42",x"00"),
  1518 => (x"20",x"20",x"20",x"54"),
  1519 => (x"4d",x"4f",x"52",x"20"),
  1520 => (x"61",x"6f",x"4c",x"00"),
  1521 => (x"2e",x"2a",x"20",x"64"),
  1522 => (x"f0",x"fe",x"1e",x"00"),
  1523 => (x"cd",x"78",x"c0",x"48"),
  1524 => (x"26",x"09",x"79",x"09"),
  1525 => (x"fe",x"1e",x"1e",x"4f"),
  1526 => (x"48",x"7e",x"bf",x"f0"),
  1527 => (x"1e",x"4f",x"26",x"26"),
  1528 => (x"c1",x"48",x"f0",x"fe"),
  1529 => (x"1e",x"4f",x"26",x"78"),
  1530 => (x"c0",x"48",x"f0",x"fe"),
  1531 => (x"1e",x"4f",x"26",x"78"),
  1532 => (x"52",x"c0",x"4a",x"71"),
  1533 => (x"0e",x"4f",x"26",x"52"),
  1534 => (x"5d",x"5c",x"5b",x"5e"),
  1535 => (x"71",x"86",x"f4",x"0e"),
  1536 => (x"7e",x"6d",x"97",x"4d"),
  1537 => (x"97",x"4c",x"a5",x"c1"),
  1538 => (x"a6",x"c8",x"48",x"6c"),
  1539 => (x"c4",x"48",x"6e",x"58"),
  1540 => (x"c5",x"05",x"a8",x"66"),
  1541 => (x"c0",x"48",x"ff",x"87"),
  1542 => (x"ca",x"ff",x"87",x"e6"),
  1543 => (x"49",x"a5",x"c2",x"87"),
  1544 => (x"71",x"4b",x"6c",x"97"),
  1545 => (x"6b",x"97",x"4b",x"a3"),
  1546 => (x"7e",x"6c",x"97",x"4b"),
  1547 => (x"80",x"c1",x"48",x"6e"),
  1548 => (x"c7",x"58",x"a6",x"c8"),
  1549 => (x"58",x"a6",x"cc",x"98"),
  1550 => (x"fe",x"7c",x"97",x"70"),
  1551 => (x"48",x"73",x"87",x"e1"),
  1552 => (x"4d",x"26",x"8e",x"f4"),
  1553 => (x"4b",x"26",x"4c",x"26"),
  1554 => (x"5e",x"0e",x"4f",x"26"),
  1555 => (x"f4",x"0e",x"5c",x"5b"),
  1556 => (x"d8",x"4c",x"71",x"86"),
  1557 => (x"ff",x"c3",x"4a",x"66"),
  1558 => (x"4b",x"a4",x"c2",x"9a"),
  1559 => (x"73",x"49",x"6c",x"97"),
  1560 => (x"51",x"72",x"49",x"a1"),
  1561 => (x"6e",x"7e",x"6c",x"97"),
  1562 => (x"c8",x"80",x"c1",x"48"),
  1563 => (x"98",x"c7",x"58",x"a6"),
  1564 => (x"70",x"58",x"a6",x"cc"),
  1565 => (x"ff",x"8e",x"f4",x"54"),
  1566 => (x"1e",x"1e",x"87",x"ca"),
  1567 => (x"e0",x"87",x"e8",x"fd"),
  1568 => (x"c0",x"49",x"4a",x"bf"),
  1569 => (x"02",x"99",x"c0",x"e0"),
  1570 => (x"1e",x"72",x"87",x"cb"),
  1571 => (x"49",x"f7",x"ec",x"c2"),
  1572 => (x"c4",x"87",x"f7",x"fe"),
  1573 => (x"87",x"fd",x"fc",x"86"),
  1574 => (x"c2",x"fd",x"7e",x"70"),
  1575 => (x"4f",x"26",x"26",x"87"),
  1576 => (x"f7",x"ec",x"c2",x"1e"),
  1577 => (x"87",x"c7",x"fd",x"49"),
  1578 => (x"49",x"fa",x"e1",x"c1"),
  1579 => (x"c5",x"87",x"da",x"fc"),
  1580 => (x"4f",x"26",x"87",x"d9"),
  1581 => (x"5c",x"5b",x"5e",x"0e"),
  1582 => (x"ed",x"c2",x"0e",x"5d"),
  1583 => (x"c1",x"4a",x"bf",x"d6"),
  1584 => (x"49",x"bf",x"c8",x"e4"),
  1585 => (x"71",x"bc",x"72",x"4c"),
  1586 => (x"87",x"db",x"fc",x"4d"),
  1587 => (x"49",x"74",x"4b",x"c0"),
  1588 => (x"d5",x"02",x"99",x"d0"),
  1589 => (x"d0",x"49",x"75",x"87"),
  1590 => (x"c0",x"1e",x"71",x"99"),
  1591 => (x"da",x"ea",x"c1",x"1e"),
  1592 => (x"12",x"82",x"73",x"4a"),
  1593 => (x"87",x"e4",x"c0",x"49"),
  1594 => (x"2c",x"c1",x"86",x"c8"),
  1595 => (x"ab",x"c8",x"83",x"2d"),
  1596 => (x"87",x"da",x"ff",x"04"),
  1597 => (x"c1",x"87",x"e8",x"fb"),
  1598 => (x"c2",x"48",x"c8",x"e4"),
  1599 => (x"78",x"bf",x"d6",x"ed"),
  1600 => (x"4c",x"26",x"4d",x"26"),
  1601 => (x"4f",x"26",x"4b",x"26"),
  1602 => (x"00",x"00",x"00",x"00"),
  1603 => (x"48",x"d0",x"ff",x"1e"),
  1604 => (x"ff",x"78",x"e1",x"c8"),
  1605 => (x"78",x"c5",x"48",x"d4"),
  1606 => (x"c3",x"02",x"66",x"c4"),
  1607 => (x"78",x"e0",x"c3",x"87"),
  1608 => (x"c6",x"02",x"66",x"c8"),
  1609 => (x"48",x"d4",x"ff",x"87"),
  1610 => (x"ff",x"78",x"f0",x"c3"),
  1611 => (x"78",x"71",x"48",x"d4"),
  1612 => (x"c8",x"48",x"d0",x"ff"),
  1613 => (x"e0",x"c0",x"78",x"e1"),
  1614 => (x"0e",x"4f",x"26",x"78"),
  1615 => (x"0e",x"5c",x"5b",x"5e"),
  1616 => (x"ec",x"c2",x"4c",x"71"),
  1617 => (x"ee",x"fa",x"49",x"f7"),
  1618 => (x"c0",x"4a",x"70",x"87"),
  1619 => (x"c2",x"04",x"aa",x"b7"),
  1620 => (x"e0",x"c3",x"87",x"e3"),
  1621 => (x"87",x"c9",x"05",x"aa"),
  1622 => (x"48",x"fe",x"e7",x"c1"),
  1623 => (x"d4",x"c2",x"78",x"c1"),
  1624 => (x"aa",x"f0",x"c3",x"87"),
  1625 => (x"c1",x"87",x"c9",x"05"),
  1626 => (x"c1",x"48",x"fa",x"e7"),
  1627 => (x"87",x"f5",x"c1",x"78"),
  1628 => (x"bf",x"fe",x"e7",x"c1"),
  1629 => (x"72",x"87",x"c7",x"02"),
  1630 => (x"b3",x"c0",x"c2",x"4b"),
  1631 => (x"4b",x"72",x"87",x"c2"),
  1632 => (x"d1",x"05",x"9c",x"74"),
  1633 => (x"fa",x"e7",x"c1",x"87"),
  1634 => (x"e7",x"c1",x"1e",x"bf"),
  1635 => (x"72",x"1e",x"bf",x"fe"),
  1636 => (x"87",x"f8",x"fd",x"49"),
  1637 => (x"e7",x"c1",x"86",x"c8"),
  1638 => (x"c0",x"02",x"bf",x"fa"),
  1639 => (x"49",x"73",x"87",x"e0"),
  1640 => (x"91",x"29",x"b7",x"c4"),
  1641 => (x"81",x"da",x"e9",x"c1"),
  1642 => (x"9a",x"cf",x"4a",x"73"),
  1643 => (x"48",x"c1",x"92",x"c2"),
  1644 => (x"4a",x"70",x"30",x"72"),
  1645 => (x"48",x"72",x"ba",x"ff"),
  1646 => (x"79",x"70",x"98",x"69"),
  1647 => (x"49",x"73",x"87",x"db"),
  1648 => (x"91",x"29",x"b7",x"c4"),
  1649 => (x"81",x"da",x"e9",x"c1"),
  1650 => (x"9a",x"cf",x"4a",x"73"),
  1651 => (x"48",x"c3",x"92",x"c2"),
  1652 => (x"4a",x"70",x"30",x"72"),
  1653 => (x"70",x"b0",x"69",x"48"),
  1654 => (x"fe",x"e7",x"c1",x"79"),
  1655 => (x"c1",x"78",x"c0",x"48"),
  1656 => (x"c0",x"48",x"fa",x"e7"),
  1657 => (x"f7",x"ec",x"c2",x"78"),
  1658 => (x"87",x"cb",x"f8",x"49"),
  1659 => (x"b7",x"c0",x"4a",x"70"),
  1660 => (x"dd",x"fd",x"03",x"aa"),
  1661 => (x"fc",x"48",x"c0",x"87"),
  1662 => (x"00",x"00",x"87",x"c8"),
  1663 => (x"00",x"00",x"00",x"00"),
  1664 => (x"71",x"1e",x"00",x"00"),
  1665 => (x"f2",x"fc",x"49",x"4a"),
  1666 => (x"1e",x"4f",x"26",x"87"),
  1667 => (x"49",x"72",x"4a",x"c0"),
  1668 => (x"e9",x"c1",x"91",x"c4"),
  1669 => (x"79",x"c0",x"81",x"da"),
  1670 => (x"b7",x"d0",x"82",x"c1"),
  1671 => (x"87",x"ee",x"04",x"aa"),
  1672 => (x"5e",x"0e",x"4f",x"26"),
  1673 => (x"0e",x"5d",x"5c",x"5b"),
  1674 => (x"fa",x"f6",x"4d",x"71"),
  1675 => (x"c4",x"4a",x"75",x"87"),
  1676 => (x"c1",x"92",x"2a",x"b7"),
  1677 => (x"75",x"82",x"da",x"e9"),
  1678 => (x"c2",x"9c",x"cf",x"4c"),
  1679 => (x"4b",x"49",x"6a",x"94"),
  1680 => (x"9b",x"c3",x"2b",x"74"),
  1681 => (x"30",x"74",x"48",x"c2"),
  1682 => (x"bc",x"ff",x"4c",x"70"),
  1683 => (x"98",x"71",x"48",x"74"),
  1684 => (x"ca",x"f6",x"7a",x"70"),
  1685 => (x"fa",x"48",x"73",x"87"),
  1686 => (x"00",x"00",x"87",x"e6"),
  1687 => (x"80",x"80",x"00",x"00"),
  1688 => (x"80",x"80",x"80",x"80"),
  1689 => (x"80",x"80",x"80",x"80"),
  1690 => (x"80",x"80",x"80",x"80"),
  1691 => (x"80",x"80",x"80",x"80"),
  1692 => (x"80",x"80",x"80",x"80"),
  1693 => (x"80",x"80",x"80",x"80"),
  1694 => (x"80",x"80",x"80",x"80"),
  1695 => (x"80",x"80",x"80",x"80"),
  1696 => (x"80",x"80",x"80",x"80"),
  1697 => (x"80",x"80",x"80",x"80"),
  1698 => (x"80",x"80",x"80",x"80"),
  1699 => (x"80",x"80",x"80",x"80"),
  1700 => (x"80",x"80",x"80",x"80"),
  1701 => (x"80",x"80",x"80",x"80"),
  1702 => (x"1e",x"16",x"80",x"80"),
  1703 => (x"36",x"2e",x"25",x"26"),
  1704 => (x"ff",x"1e",x"3e",x"3d"),
  1705 => (x"e1",x"c8",x"48",x"d0"),
  1706 => (x"ff",x"48",x"71",x"78"),
  1707 => (x"26",x"78",x"08",x"d4"),
  1708 => (x"d0",x"ff",x"1e",x"4f"),
  1709 => (x"78",x"e1",x"c8",x"48"),
  1710 => (x"d4",x"ff",x"48",x"71"),
  1711 => (x"66",x"c4",x"78",x"08"),
  1712 => (x"08",x"d4",x"ff",x"48"),
  1713 => (x"1e",x"4f",x"26",x"78"),
  1714 => (x"66",x"c4",x"4a",x"71"),
  1715 => (x"49",x"72",x"1e",x"49"),
  1716 => (x"ff",x"87",x"de",x"ff"),
  1717 => (x"e0",x"c0",x"48",x"d0"),
  1718 => (x"4f",x"26",x"26",x"78"),
  1719 => (x"c2",x"4a",x"71",x"1e"),
  1720 => (x"c3",x"03",x"aa",x"b7"),
  1721 => (x"87",x"c2",x"82",x"87"),
  1722 => (x"66",x"c4",x"82",x"ce"),
  1723 => (x"ff",x"49",x"72",x"1e"),
  1724 => (x"26",x"26",x"87",x"d5"),
  1725 => (x"d4",x"ff",x"1e",x"4f"),
  1726 => (x"7a",x"ff",x"c3",x"4a"),
  1727 => (x"c8",x"48",x"d0",x"ff"),
  1728 => (x"7a",x"de",x"78",x"e1"),
  1729 => (x"bf",x"c1",x"ed",x"c2"),
  1730 => (x"c8",x"48",x"49",x"7a"),
  1731 => (x"71",x"7a",x"70",x"28"),
  1732 => (x"70",x"28",x"d0",x"48"),
  1733 => (x"d8",x"48",x"71",x"7a"),
  1734 => (x"ff",x"7a",x"70",x"28"),
  1735 => (x"e0",x"c0",x"48",x"d0"),
  1736 => (x"0e",x"4f",x"26",x"78"),
  1737 => (x"5d",x"5c",x"5b",x"5e"),
  1738 => (x"c2",x"4c",x"71",x"0e"),
  1739 => (x"4d",x"bf",x"c1",x"ed"),
  1740 => (x"d0",x"2b",x"74",x"4b"),
  1741 => (x"83",x"c1",x"9b",x"66"),
  1742 => (x"04",x"ab",x"66",x"d4"),
  1743 => (x"4b",x"c0",x"87",x"c2"),
  1744 => (x"66",x"d0",x"4a",x"74"),
  1745 => (x"ff",x"31",x"72",x"49"),
  1746 => (x"73",x"99",x"75",x"b9"),
  1747 => (x"70",x"30",x"72",x"48"),
  1748 => (x"b0",x"71",x"48",x"4a"),
  1749 => (x"58",x"c5",x"ed",x"c2"),
  1750 => (x"26",x"87",x"da",x"fe"),
  1751 => (x"26",x"4c",x"26",x"4d"),
  1752 => (x"1e",x"4f",x"26",x"4b"),
  1753 => (x"c8",x"48",x"d0",x"ff"),
  1754 => (x"48",x"71",x"78",x"c9"),
  1755 => (x"78",x"08",x"d4",x"ff"),
  1756 => (x"71",x"1e",x"4f",x"26"),
  1757 => (x"87",x"eb",x"49",x"4a"),
  1758 => (x"c8",x"48",x"d0",x"ff"),
  1759 => (x"1e",x"4f",x"26",x"78"),
  1760 => (x"4b",x"71",x"1e",x"73"),
  1761 => (x"bf",x"d1",x"ed",x"c2"),
  1762 => (x"c2",x"87",x"c3",x"02"),
  1763 => (x"d0",x"ff",x"87",x"eb"),
  1764 => (x"78",x"c9",x"c8",x"48"),
  1765 => (x"e0",x"c0",x"49",x"73"),
  1766 => (x"48",x"d4",x"ff",x"b1"),
  1767 => (x"ed",x"c2",x"78",x"71"),
  1768 => (x"78",x"c0",x"48",x"c5"),
  1769 => (x"c5",x"02",x"66",x"c8"),
  1770 => (x"49",x"ff",x"c3",x"87"),
  1771 => (x"49",x"c0",x"87",x"c2"),
  1772 => (x"59",x"cd",x"ed",x"c2"),
  1773 => (x"c6",x"02",x"66",x"cc"),
  1774 => (x"d5",x"d5",x"c5",x"87"),
  1775 => (x"cf",x"87",x"c4",x"4a"),
  1776 => (x"c2",x"4a",x"ff",x"ff"),
  1777 => (x"c2",x"5a",x"d1",x"ed"),
  1778 => (x"c1",x"48",x"d1",x"ed"),
  1779 => (x"26",x"87",x"c4",x"78"),
  1780 => (x"26",x"4c",x"26",x"4d"),
  1781 => (x"0e",x"4f",x"26",x"4b"),
  1782 => (x"5d",x"5c",x"5b",x"5e"),
  1783 => (x"c2",x"4a",x"71",x"0e"),
  1784 => (x"4c",x"bf",x"cd",x"ed"),
  1785 => (x"cb",x"02",x"9a",x"72"),
  1786 => (x"91",x"c8",x"49",x"87"),
  1787 => (x"4b",x"f5",x"ed",x"c1"),
  1788 => (x"87",x"c4",x"83",x"71"),
  1789 => (x"4b",x"f5",x"f1",x"c1"),
  1790 => (x"49",x"13",x"4d",x"c0"),
  1791 => (x"ed",x"c2",x"99",x"74"),
  1792 => (x"ff",x"b9",x"bf",x"c9"),
  1793 => (x"78",x"71",x"48",x"d4"),
  1794 => (x"85",x"2c",x"b7",x"c1"),
  1795 => (x"04",x"ad",x"b7",x"c8"),
  1796 => (x"ed",x"c2",x"87",x"e8"),
  1797 => (x"c8",x"48",x"bf",x"c5"),
  1798 => (x"c9",x"ed",x"c2",x"80"),
  1799 => (x"87",x"ef",x"fe",x"58"),
  1800 => (x"71",x"1e",x"73",x"1e"),
  1801 => (x"9a",x"4a",x"13",x"4b"),
  1802 => (x"72",x"87",x"cb",x"02"),
  1803 => (x"87",x"e7",x"fe",x"49"),
  1804 => (x"05",x"9a",x"4a",x"13"),
  1805 => (x"da",x"fe",x"87",x"f5"),
  1806 => (x"ed",x"c2",x"1e",x"87"),
  1807 => (x"c2",x"49",x"bf",x"c5"),
  1808 => (x"c1",x"48",x"c5",x"ed"),
  1809 => (x"c0",x"c4",x"78",x"a1"),
  1810 => (x"db",x"03",x"a9",x"b7"),
  1811 => (x"48",x"d4",x"ff",x"87"),
  1812 => (x"bf",x"c9",x"ed",x"c2"),
  1813 => (x"c5",x"ed",x"c2",x"78"),
  1814 => (x"ed",x"c2",x"49",x"bf"),
  1815 => (x"a1",x"c1",x"48",x"c5"),
  1816 => (x"b7",x"c0",x"c4",x"78"),
  1817 => (x"87",x"e5",x"04",x"a9"),
  1818 => (x"c8",x"48",x"d0",x"ff"),
  1819 => (x"d1",x"ed",x"c2",x"78"),
  1820 => (x"26",x"78",x"c0",x"48"),
  1821 => (x"00",x"00",x"00",x"4f"),
  1822 => (x"00",x"00",x"00",x"00"),
  1823 => (x"00",x"00",x"00",x"00"),
  1824 => (x"00",x"00",x"5f",x"5f"),
  1825 => (x"03",x"03",x"00",x"00"),
  1826 => (x"00",x"03",x"03",x"00"),
  1827 => (x"7f",x"7f",x"14",x"00"),
  1828 => (x"14",x"7f",x"7f",x"14"),
  1829 => (x"2e",x"24",x"00",x"00"),
  1830 => (x"12",x"3a",x"6b",x"6b"),
  1831 => (x"36",x"6a",x"4c",x"00"),
  1832 => (x"32",x"56",x"6c",x"18"),
  1833 => (x"4f",x"7e",x"30",x"00"),
  1834 => (x"68",x"3a",x"77",x"59"),
  1835 => (x"04",x"00",x"00",x"40"),
  1836 => (x"00",x"00",x"03",x"07"),
  1837 => (x"1c",x"00",x"00",x"00"),
  1838 => (x"00",x"41",x"63",x"3e"),
  1839 => (x"41",x"00",x"00",x"00"),
  1840 => (x"00",x"1c",x"3e",x"63"),
  1841 => (x"3e",x"2a",x"08",x"00"),
  1842 => (x"2a",x"3e",x"1c",x"1c"),
  1843 => (x"08",x"08",x"00",x"08"),
  1844 => (x"08",x"08",x"3e",x"3e"),
  1845 => (x"80",x"00",x"00",x"00"),
  1846 => (x"00",x"00",x"60",x"e0"),
  1847 => (x"08",x"08",x"00",x"00"),
  1848 => (x"08",x"08",x"08",x"08"),
  1849 => (x"00",x"00",x"00",x"00"),
  1850 => (x"00",x"00",x"60",x"60"),
  1851 => (x"30",x"60",x"40",x"00"),
  1852 => (x"03",x"06",x"0c",x"18"),
  1853 => (x"7f",x"3e",x"00",x"01"),
  1854 => (x"3e",x"7f",x"4d",x"59"),
  1855 => (x"06",x"04",x"00",x"00"),
  1856 => (x"00",x"00",x"7f",x"7f"),
  1857 => (x"63",x"42",x"00",x"00"),
  1858 => (x"46",x"4f",x"59",x"71"),
  1859 => (x"63",x"22",x"00",x"00"),
  1860 => (x"36",x"7f",x"49",x"49"),
  1861 => (x"16",x"1c",x"18",x"00"),
  1862 => (x"10",x"7f",x"7f",x"13"),
  1863 => (x"67",x"27",x"00",x"00"),
  1864 => (x"39",x"7d",x"45",x"45"),
  1865 => (x"7e",x"3c",x"00",x"00"),
  1866 => (x"30",x"79",x"49",x"4b"),
  1867 => (x"01",x"01",x"00",x"00"),
  1868 => (x"07",x"0f",x"79",x"71"),
  1869 => (x"7f",x"36",x"00",x"00"),
  1870 => (x"36",x"7f",x"49",x"49"),
  1871 => (x"4f",x"06",x"00",x"00"),
  1872 => (x"1e",x"3f",x"69",x"49"),
  1873 => (x"00",x"00",x"00",x"00"),
  1874 => (x"00",x"00",x"66",x"66"),
  1875 => (x"80",x"00",x"00",x"00"),
  1876 => (x"00",x"00",x"66",x"e6"),
  1877 => (x"08",x"08",x"00",x"00"),
  1878 => (x"22",x"22",x"14",x"14"),
  1879 => (x"14",x"14",x"00",x"00"),
  1880 => (x"14",x"14",x"14",x"14"),
  1881 => (x"22",x"22",x"00",x"00"),
  1882 => (x"08",x"08",x"14",x"14"),
  1883 => (x"03",x"02",x"00",x"00"),
  1884 => (x"06",x"0f",x"59",x"51"),
  1885 => (x"41",x"7f",x"3e",x"00"),
  1886 => (x"1e",x"1f",x"55",x"5d"),
  1887 => (x"7f",x"7e",x"00",x"00"),
  1888 => (x"7e",x"7f",x"09",x"09"),
  1889 => (x"7f",x"7f",x"00",x"00"),
  1890 => (x"36",x"7f",x"49",x"49"),
  1891 => (x"3e",x"1c",x"00",x"00"),
  1892 => (x"41",x"41",x"41",x"63"),
  1893 => (x"7f",x"7f",x"00",x"00"),
  1894 => (x"1c",x"3e",x"63",x"41"),
  1895 => (x"7f",x"7f",x"00",x"00"),
  1896 => (x"41",x"41",x"49",x"49"),
  1897 => (x"7f",x"7f",x"00",x"00"),
  1898 => (x"01",x"01",x"09",x"09"),
  1899 => (x"7f",x"3e",x"00",x"00"),
  1900 => (x"7a",x"7b",x"49",x"41"),
  1901 => (x"7f",x"7f",x"00",x"00"),
  1902 => (x"7f",x"7f",x"08",x"08"),
  1903 => (x"41",x"00",x"00",x"00"),
  1904 => (x"00",x"41",x"7f",x"7f"),
  1905 => (x"60",x"20",x"00",x"00"),
  1906 => (x"3f",x"7f",x"40",x"40"),
  1907 => (x"08",x"7f",x"7f",x"00"),
  1908 => (x"41",x"63",x"36",x"1c"),
  1909 => (x"7f",x"7f",x"00",x"00"),
  1910 => (x"40",x"40",x"40",x"40"),
  1911 => (x"06",x"7f",x"7f",x"00"),
  1912 => (x"7f",x"7f",x"06",x"0c"),
  1913 => (x"06",x"7f",x"7f",x"00"),
  1914 => (x"7f",x"7f",x"18",x"0c"),
  1915 => (x"7f",x"3e",x"00",x"00"),
  1916 => (x"3e",x"7f",x"41",x"41"),
  1917 => (x"7f",x"7f",x"00",x"00"),
  1918 => (x"06",x"0f",x"09",x"09"),
  1919 => (x"41",x"7f",x"3e",x"00"),
  1920 => (x"40",x"7e",x"7f",x"61"),
  1921 => (x"7f",x"7f",x"00",x"00"),
  1922 => (x"66",x"7f",x"19",x"09"),
  1923 => (x"6f",x"26",x"00",x"00"),
  1924 => (x"32",x"7b",x"59",x"4d"),
  1925 => (x"01",x"01",x"00",x"00"),
  1926 => (x"01",x"01",x"7f",x"7f"),
  1927 => (x"7f",x"3f",x"00",x"00"),
  1928 => (x"3f",x"7f",x"40",x"40"),
  1929 => (x"3f",x"0f",x"00",x"00"),
  1930 => (x"0f",x"3f",x"70",x"70"),
  1931 => (x"30",x"7f",x"7f",x"00"),
  1932 => (x"7f",x"7f",x"30",x"18"),
  1933 => (x"36",x"63",x"41",x"00"),
  1934 => (x"63",x"36",x"1c",x"1c"),
  1935 => (x"06",x"03",x"01",x"41"),
  1936 => (x"03",x"06",x"7c",x"7c"),
  1937 => (x"59",x"71",x"61",x"01"),
  1938 => (x"41",x"43",x"47",x"4d"),
  1939 => (x"7f",x"00",x"00",x"00"),
  1940 => (x"00",x"41",x"41",x"7f"),
  1941 => (x"06",x"03",x"01",x"00"),
  1942 => (x"60",x"30",x"18",x"0c"),
  1943 => (x"41",x"00",x"00",x"40"),
  1944 => (x"00",x"7f",x"7f",x"41"),
  1945 => (x"06",x"0c",x"08",x"00"),
  1946 => (x"08",x"0c",x"06",x"03"),
  1947 => (x"80",x"80",x"80",x"00"),
  1948 => (x"80",x"80",x"80",x"80"),
  1949 => (x"00",x"00",x"00",x"00"),
  1950 => (x"00",x"04",x"07",x"03"),
  1951 => (x"74",x"20",x"00",x"00"),
  1952 => (x"78",x"7c",x"54",x"54"),
  1953 => (x"7f",x"7f",x"00",x"00"),
  1954 => (x"38",x"7c",x"44",x"44"),
  1955 => (x"7c",x"38",x"00",x"00"),
  1956 => (x"00",x"44",x"44",x"44"),
  1957 => (x"7c",x"38",x"00",x"00"),
  1958 => (x"7f",x"7f",x"44",x"44"),
  1959 => (x"7c",x"38",x"00",x"00"),
  1960 => (x"18",x"5c",x"54",x"54"),
  1961 => (x"7e",x"04",x"00",x"00"),
  1962 => (x"00",x"05",x"05",x"7f"),
  1963 => (x"bc",x"18",x"00",x"00"),
  1964 => (x"7c",x"fc",x"a4",x"a4"),
  1965 => (x"7f",x"7f",x"00",x"00"),
  1966 => (x"78",x"7c",x"04",x"04"),
  1967 => (x"00",x"00",x"00",x"00"),
  1968 => (x"00",x"40",x"7d",x"3d"),
  1969 => (x"80",x"80",x"00",x"00"),
  1970 => (x"00",x"7d",x"fd",x"80"),
  1971 => (x"7f",x"7f",x"00",x"00"),
  1972 => (x"44",x"6c",x"38",x"10"),
  1973 => (x"00",x"00",x"00",x"00"),
  1974 => (x"00",x"40",x"7f",x"3f"),
  1975 => (x"0c",x"7c",x"7c",x"00"),
  1976 => (x"78",x"7c",x"0c",x"18"),
  1977 => (x"7c",x"7c",x"00",x"00"),
  1978 => (x"78",x"7c",x"04",x"04"),
  1979 => (x"7c",x"38",x"00",x"00"),
  1980 => (x"38",x"7c",x"44",x"44"),
  1981 => (x"fc",x"fc",x"00",x"00"),
  1982 => (x"18",x"3c",x"24",x"24"),
  1983 => (x"3c",x"18",x"00",x"00"),
  1984 => (x"fc",x"fc",x"24",x"24"),
  1985 => (x"7c",x"7c",x"00",x"00"),
  1986 => (x"08",x"0c",x"04",x"04"),
  1987 => (x"5c",x"48",x"00",x"00"),
  1988 => (x"20",x"74",x"54",x"54"),
  1989 => (x"3f",x"04",x"00",x"00"),
  1990 => (x"00",x"44",x"44",x"7f"),
  1991 => (x"7c",x"3c",x"00",x"00"),
  1992 => (x"7c",x"7c",x"40",x"40"),
  1993 => (x"3c",x"1c",x"00",x"00"),
  1994 => (x"1c",x"3c",x"60",x"60"),
  1995 => (x"60",x"7c",x"3c",x"00"),
  1996 => (x"3c",x"7c",x"60",x"30"),
  1997 => (x"38",x"6c",x"44",x"00"),
  1998 => (x"44",x"6c",x"38",x"10"),
  1999 => (x"bc",x"1c",x"00",x"00"),
  2000 => (x"1c",x"3c",x"60",x"e0"),
  2001 => (x"64",x"44",x"00",x"00"),
  2002 => (x"44",x"4c",x"5c",x"74"),
  2003 => (x"08",x"08",x"00",x"00"),
  2004 => (x"41",x"41",x"77",x"3e"),
  2005 => (x"00",x"00",x"00",x"00"),
  2006 => (x"00",x"00",x"7f",x"7f"),
  2007 => (x"41",x"41",x"00",x"00"),
  2008 => (x"08",x"08",x"3e",x"77"),
  2009 => (x"01",x"01",x"02",x"00"),
  2010 => (x"01",x"02",x"02",x"03"),
  2011 => (x"7f",x"7f",x"7f",x"00"),
  2012 => (x"7f",x"7f",x"7f",x"7f"),
  2013 => (x"1c",x"08",x"08",x"00"),
  2014 => (x"7f",x"3e",x"3e",x"1c"),
  2015 => (x"3e",x"7f",x"7f",x"7f"),
  2016 => (x"08",x"1c",x"1c",x"3e"),
  2017 => (x"18",x"10",x"00",x"08"),
  2018 => (x"10",x"18",x"7c",x"7c"),
  2019 => (x"30",x"10",x"00",x"00"),
  2020 => (x"10",x"30",x"7c",x"7c"),
  2021 => (x"60",x"30",x"10",x"00"),
  2022 => (x"06",x"1e",x"78",x"60"),
  2023 => (x"3c",x"66",x"42",x"00"),
  2024 => (x"42",x"66",x"3c",x"18"),
  2025 => (x"6a",x"38",x"78",x"00"),
  2026 => (x"38",x"6c",x"c6",x"c2"),
  2027 => (x"00",x"00",x"60",x"00"),
  2028 => (x"60",x"00",x"00",x"60"),
  2029 => (x"5b",x"5e",x"0e",x"00"),
  2030 => (x"1e",x"0e",x"5d",x"5c"),
  2031 => (x"ed",x"c2",x"4c",x"71"),
  2032 => (x"c0",x"4d",x"bf",x"e2"),
  2033 => (x"74",x"1e",x"c0",x"4b"),
  2034 => (x"87",x"c7",x"02",x"ab"),
  2035 => (x"c0",x"48",x"a6",x"c4"),
  2036 => (x"c4",x"87",x"c5",x"78"),
  2037 => (x"78",x"c1",x"48",x"a6"),
  2038 => (x"73",x"1e",x"66",x"c4"),
  2039 => (x"87",x"df",x"ee",x"49"),
  2040 => (x"e0",x"c0",x"86",x"c8"),
  2041 => (x"87",x"ef",x"ef",x"49"),
  2042 => (x"6a",x"4a",x"a5",x"c4"),
  2043 => (x"87",x"f0",x"f0",x"49"),
  2044 => (x"cb",x"87",x"c6",x"f1"),
  2045 => (x"c8",x"83",x"c1",x"85"),
  2046 => (x"ff",x"04",x"ab",x"b7"),
  2047 => (x"26",x"26",x"87",x"c7"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

