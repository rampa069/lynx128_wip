library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom1 is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom1 is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0487da01",
     1 => x"580e87dd",
     2 => x"0e5a595e",
     3 => x"00002927",
     4 => x"4a260f00",
     5 => x"48264926",
     6 => x"082680ff",
     7 => x"002d274f",
     8 => x"274f0000",
     9 => x"0000002a",
    10 => x"fd004f4f",
    11 => x"d4eec287",
    12 => x"86c0c64e",
    13 => x"49d4eec2",
    14 => x"48f4dbc2",
    15 => x"4040c089",
    16 => x"89d04040",
    17 => x"c187f603",
    18 => x"0087dfdb",
    19 => x"1e87fc98",
    20 => x"1e731e72",
    21 => x"02114812",
    22 => x"c34b87ca",
    23 => x"739b98df",
    24 => x"87f00288",
    25 => x"4a264b26",
    26 => x"731e4f26",
    27 => x"c11e721e",
    28 => x"87ca048b",
    29 => x"02114812",
    30 => x"028887c4",
    31 => x"4a2687f1",
    32 => x"4f264b26",
    33 => x"731e741e",
    34 => x"c11e721e",
    35 => x"87d0048b",
    36 => x"02114812",
    37 => x"c34c87ca",
    38 => x"749c98df",
    39 => x"87eb0288",
    40 => x"4b264a26",
    41 => x"4f264c26",
    42 => x"8148731e",
    43 => x"c502a973",
    44 => x"05531287",
    45 => x"4f2687f6",
    46 => x"4a66c41e",
    47 => x"51124871",
    48 => x"2687fb05",
    49 => x"66c41e4f",
    50 => x"ff48114a",
    51 => x"c17808d4",
    52 => x"87f5058a",
    53 => x"c41e4f26",
    54 => x"d4ff4a66",
    55 => x"78ffc348",
    56 => x"8ac15168",
    57 => x"2687f305",
    58 => x"1e731e4f",
    59 => x"c34bd4ff",
    60 => x"4a6b7bff",
    61 => x"6b7bffc3",
    62 => x"7232c849",
    63 => x"7bffc3b1",
    64 => x"31c84a6b",
    65 => x"ffc3b271",
    66 => x"c8496b7b",
    67 => x"71b17232",
    68 => x"2687c448",
    69 => x"264c264d",
    70 => x"0e4f264b",
    71 => x"5d5c5b5e",
    72 => x"ff4a710e",
    73 => x"49724cd4",
    74 => x"7199ffc3",
    75 => x"f4dbc27c",
    76 => x"87c805bf",
    77 => x"c94866d0",
    78 => x"58a6d430",
    79 => x"d84966d0",
    80 => x"99ffc329",
    81 => x"66d07c71",
    82 => x"c329d049",
    83 => x"7c7199ff",
    84 => x"c84966d0",
    85 => x"99ffc329",
    86 => x"66d07c71",
    87 => x"99ffc349",
    88 => x"49727c71",
    89 => x"ffc329d0",
    90 => x"6c7c7199",
    91 => x"fff0c94b",
    92 => x"abffc34d",
    93 => x"c387d005",
    94 => x"4b6c7cff",
    95 => x"c6028dc1",
    96 => x"abffc387",
    97 => x"7387f002",
    98 => x"87c7fe48",
    99 => x"ff49c01e",
   100 => x"ffc348d4",
   101 => x"c381c178",
   102 => x"04a9b7c8",
   103 => x"4f2687f1",
   104 => x"e71e731e",
   105 => x"dff8c487",
   106 => x"c01ec04b",
   107 => x"f7c1f0ff",
   108 => x"87e7fd49",
   109 => x"a8c186c4",
   110 => x"87eac005",
   111 => x"c348d4ff",
   112 => x"c0c178ff",
   113 => x"c0c0c0c0",
   114 => x"f0e1c01e",
   115 => x"fd49e9c1",
   116 => x"86c487c9",
   117 => x"ca059870",
   118 => x"48d4ff87",
   119 => x"c178ffc3",
   120 => x"fe87cb48",
   121 => x"8bc187e6",
   122 => x"87fdfe05",
   123 => x"e6fc48c0",
   124 => x"1e731e87",
   125 => x"c348d4ff",
   126 => x"4bd378ff",
   127 => x"ffc01ec0",
   128 => x"49c1c1f0",
   129 => x"c487d4fc",
   130 => x"05987086",
   131 => x"d4ff87ca",
   132 => x"78ffc348",
   133 => x"87cb48c1",
   134 => x"c187f1fd",
   135 => x"dbff058b",
   136 => x"fb48c087",
   137 => x"5e0e87f1",
   138 => x"ff0e5c5b",
   139 => x"dbfd4cd4",
   140 => x"1eeac687",
   141 => x"c1f0e1c0",
   142 => x"defb49c8",
   143 => x"c186c487",
   144 => x"87c802a8",
   145 => x"c087eafe",
   146 => x"87e2c148",
   147 => x"7087dafa",
   148 => x"ffffcf49",
   149 => x"a9eac699",
   150 => x"fe87c802",
   151 => x"48c087d3",
   152 => x"c387cbc1",
   153 => x"f1c07cff",
   154 => x"87f4fc4b",
   155 => x"c0029870",
   156 => x"1ec087eb",
   157 => x"c1f0ffc0",
   158 => x"defa49fa",
   159 => x"7086c487",
   160 => x"87d90598",
   161 => x"6c7cffc3",
   162 => x"7cffc349",
   163 => x"c17c7c7c",
   164 => x"c40299c0",
   165 => x"d548c187",
   166 => x"d148c087",
   167 => x"05abc287",
   168 => x"48c087c4",
   169 => x"8bc187c8",
   170 => x"87fdfe05",
   171 => x"e4f948c0",
   172 => x"1e731e87",
   173 => x"48f4dbc2",
   174 => x"4bc778c1",
   175 => x"c248d0ff",
   176 => x"87c8fb78",
   177 => x"c348d0ff",
   178 => x"c01ec078",
   179 => x"c0c1d0e5",
   180 => x"87c7f949",
   181 => x"a8c186c4",
   182 => x"4b87c105",
   183 => x"c505abc2",
   184 => x"c048c087",
   185 => x"8bc187f9",
   186 => x"87d0ff05",
   187 => x"c287f7fc",
   188 => x"7058f8db",
   189 => x"87cd0598",
   190 => x"ffc01ec1",
   191 => x"49d0c1f0",
   192 => x"c487d8f8",
   193 => x"48d4ff86",
   194 => x"c478ffc3",
   195 => x"dbc287e0",
   196 => x"d0ff58fc",
   197 => x"ff78c248",
   198 => x"ffc348d4",
   199 => x"f748c178",
   200 => x"5e0e87f5",
   201 => x"0e5d5c5b",
   202 => x"ffc34a71",
   203 => x"4cd4ff4d",
   204 => x"d0ff7c75",
   205 => x"78c3c448",
   206 => x"1e727c75",
   207 => x"c1f0ffc0",
   208 => x"d6f749d8",
   209 => x"7086c487",
   210 => x"87c50298",
   211 => x"f0c048c0",
   212 => x"c37c7587",
   213 => x"c0c87cfe",
   214 => x"4966d41e",
   215 => x"c487e6f5",
   216 => x"757c7586",
   217 => x"d87c757c",
   218 => x"754be0da",
   219 => x"99496c7c",
   220 => x"c187c505",
   221 => x"87f3058b",
   222 => x"d0ff7c75",
   223 => x"c178c248",
   224 => x"87cff648",
   225 => x"4ad4ff1e",
   226 => x"c448d0ff",
   227 => x"ffc378d1",
   228 => x"0589c17a",
   229 => x"4f2687f8",
   230 => x"711e731e",
   231 => x"cdeec54b",
   232 => x"d4ff4adf",
   233 => x"78ffc348",
   234 => x"fec34868",
   235 => x"87c502a8",
   236 => x"ed058ac1",
   237 => x"059a7287",
   238 => x"48c087c5",
   239 => x"7387eac0",
   240 => x"87cc029b",
   241 => x"731e66c8",
   242 => x"87caf449",
   243 => x"87c686c4",
   244 => x"fe4966c8",
   245 => x"d4ff87ee",
   246 => x"78ffc348",
   247 => x"059b7378",
   248 => x"d0ff87c5",
   249 => x"c178d048",
   250 => x"87ebf448",
   251 => x"711e731e",
   252 => x"ff4bc04a",
   253 => x"ffc348d4",
   254 => x"48d0ff78",
   255 => x"ff78c3c4",
   256 => x"ffc348d4",
   257 => x"c01e7278",
   258 => x"d1c1f0ff",
   259 => x"87cbf449",
   260 => x"987086c4",
   261 => x"c887cd05",
   262 => x"66cc1ec0",
   263 => x"87f8fd49",
   264 => x"4b7086c4",
   265 => x"c248d0ff",
   266 => x"f3487378",
   267 => x"5e0e87e9",
   268 => x"0e5d5c5b",
   269 => x"ffc01ec0",
   270 => x"49c9c1f0",
   271 => x"d287dcf3",
   272 => x"fcdbc21e",
   273 => x"87d0fd49",
   274 => x"4cc086c8",
   275 => x"b7d284c1",
   276 => x"87f804ac",
   277 => x"97fcdbc2",
   278 => x"c0c349bf",
   279 => x"a9c0c199",
   280 => x"87e7c005",
   281 => x"97c3dcc2",
   282 => x"31d049bf",
   283 => x"97c4dcc2",
   284 => x"32c84abf",
   285 => x"dcc2b172",
   286 => x"4abf97c5",
   287 => x"cf4c71b1",
   288 => x"9cffffff",
   289 => x"34ca84c1",
   290 => x"c287e7c1",
   291 => x"bf97c5dc",
   292 => x"c631c149",
   293 => x"c6dcc299",
   294 => x"c74abf97",
   295 => x"b1722ab7",
   296 => x"97c1dcc2",
   297 => x"cf4d4abf",
   298 => x"c2dcc29d",
   299 => x"c34abf97",
   300 => x"c232ca9a",
   301 => x"bf97c3dc",
   302 => x"7333c24b",
   303 => x"c4dcc2b2",
   304 => x"c34bbf97",
   305 => x"b7c69bc0",
   306 => x"c2b2732b",
   307 => x"7148c181",
   308 => x"c1497030",
   309 => x"70307548",
   310 => x"c14c724d",
   311 => x"c8947184",
   312 => x"06adb7c0",
   313 => x"34c187cc",
   314 => x"c0c82db7",
   315 => x"ff01adb7",
   316 => x"487487f4",
   317 => x"0e87dcf0",
   318 => x"5d5c5b5e",
   319 => x"c286f80e",
   320 => x"c048e2e4",
   321 => x"dadcc278",
   322 => x"fb49c01e",
   323 => x"86c487de",
   324 => x"c5059870",
   325 => x"c948c087",
   326 => x"4dc087ce",
   327 => x"f2c07ec1",
   328 => x"c249bfc1",
   329 => x"714ad0dd",
   330 => x"fdec4bc8",
   331 => x"05987087",
   332 => x"7ec087c2",
   333 => x"bffdf1c0",
   334 => x"ecddc249",
   335 => x"4bc8714a",
   336 => x"7087e7ec",
   337 => x"87c20598",
   338 => x"026e7ec0",
   339 => x"c287fdc0",
   340 => x"4dbfe0e3",
   341 => x"9fd8e4c2",
   342 => x"c5487ebf",
   343 => x"05a8ead6",
   344 => x"e3c287c7",
   345 => x"ce4dbfe0",
   346 => x"ca486e87",
   347 => x"02a8d5e9",
   348 => x"48c087c5",
   349 => x"c287f1c7",
   350 => x"751edadc",
   351 => x"87ecf949",
   352 => x"987086c4",
   353 => x"c087c505",
   354 => x"87dcc748",
   355 => x"bffdf1c0",
   356 => x"ecddc249",
   357 => x"4bc8714a",
   358 => x"7087cfeb",
   359 => x"87c80598",
   360 => x"48e2e4c2",
   361 => x"87da78c1",
   362 => x"bfc1f2c0",
   363 => x"d0ddc249",
   364 => x"4bc8714a",
   365 => x"7087f3ea",
   366 => x"c5c00298",
   367 => x"c648c087",
   368 => x"e4c287e6",
   369 => x"49bf97d8",
   370 => x"05a9d5c1",
   371 => x"c287cdc0",
   372 => x"bf97d9e4",
   373 => x"a9eac249",
   374 => x"87c5c002",
   375 => x"c7c648c0",
   376 => x"dadcc287",
   377 => x"487ebf97",
   378 => x"02a8e9c3",
   379 => x"6e87cec0",
   380 => x"a8ebc348",
   381 => x"87c5c002",
   382 => x"ebc548c0",
   383 => x"e5dcc287",
   384 => x"9949bf97",
   385 => x"87ccc005",
   386 => x"97e6dcc2",
   387 => x"a9c249bf",
   388 => x"87c5c002",
   389 => x"cfc548c0",
   390 => x"e7dcc287",
   391 => x"c248bf97",
   392 => x"7058dee4",
   393 => x"88c1484c",
   394 => x"58e2e4c2",
   395 => x"97e8dcc2",
   396 => x"817549bf",
   397 => x"97e9dcc2",
   398 => x"32c84abf",
   399 => x"c27ea172",
   400 => x"6e48efe8",
   401 => x"eadcc278",
   402 => x"c848bf97",
   403 => x"e4c258a6",
   404 => x"c202bfe2",
   405 => x"f1c087d4",
   406 => x"c249bffd",
   407 => x"714aecdd",
   408 => x"c5e84bc8",
   409 => x"02987087",
   410 => x"c087c5c0",
   411 => x"87f8c348",
   412 => x"bfdae4c2",
   413 => x"c3e9c24c",
   414 => x"ffdcc25c",
   415 => x"c849bf97",
   416 => x"fedcc231",
   417 => x"a14abf97",
   418 => x"c0ddc249",
   419 => x"d04abf97",
   420 => x"49a17232",
   421 => x"97c1ddc2",
   422 => x"32d84abf",
   423 => x"c449a172",
   424 => x"e8c29166",
   425 => x"c281bfef",
   426 => x"c259f7e8",
   427 => x"bf97c7dd",
   428 => x"c232c84a",
   429 => x"bf97c6dd",
   430 => x"c24aa24b",
   431 => x"bf97c8dd",
   432 => x"7333d04b",
   433 => x"ddc24aa2",
   434 => x"4bbf97c9",
   435 => x"33d89bcf",
   436 => x"c24aa273",
   437 => x"c25afbe8",
   438 => x"4abff7e8",
   439 => x"92748ac2",
   440 => x"48fbe8c2",
   441 => x"c178a172",
   442 => x"dcc287ca",
   443 => x"49bf97ec",
   444 => x"dcc231c8",
   445 => x"4abf97eb",
   446 => x"e4c249a1",
   447 => x"e4c259ea",
   448 => x"c549bfe6",
   449 => x"81ffc731",
   450 => x"e9c229c9",
   451 => x"dcc259c3",
   452 => x"4abf97f1",
   453 => x"dcc232c8",
   454 => x"4bbf97f0",
   455 => x"66c44aa2",
   456 => x"c2826e92",
   457 => x"c25affe8",
   458 => x"c048f7e8",
   459 => x"f3e8c278",
   460 => x"78a17248",
   461 => x"48c3e9c2",
   462 => x"bff7e8c2",
   463 => x"c7e9c278",
   464 => x"fbe8c248",
   465 => x"e4c278bf",
   466 => x"c002bfe2",
   467 => x"487487c9",
   468 => x"7e7030c4",
   469 => x"c287c9c0",
   470 => x"48bfffe8",
   471 => x"7e7030c4",
   472 => x"48e6e4c2",
   473 => x"48c1786e",
   474 => x"4d268ef8",
   475 => x"4b264c26",
   476 => x"5e0e4f26",
   477 => x"0e5d5c5b",
   478 => x"e4c24a71",
   479 => x"cb02bfe2",
   480 => x"c74b7287",
   481 => x"c14c722b",
   482 => x"87c99cff",
   483 => x"2bc84b72",
   484 => x"ffc34c72",
   485 => x"efe8c29c",
   486 => x"f1c083bf",
   487 => x"02abbff9",
   488 => x"f1c087d9",
   489 => x"dcc25bfd",
   490 => x"49731eda",
   491 => x"c487fdf0",
   492 => x"05987086",
   493 => x"48c087c5",
   494 => x"c287e6c0",
   495 => x"02bfe2e4",
   496 => x"497487d2",
   497 => x"dcc291c4",
   498 => x"4d6981da",
   499 => x"ffffffcf",
   500 => x"87cb9dff",
   501 => x"91c24974",
   502 => x"81dadcc2",
   503 => x"754d699f",
   504 => x"87c6fe48",
   505 => x"5c5b5e0e",
   506 => x"711e0e5d",
   507 => x"c11ec04d",
   508 => x"87eeca49",
   509 => x"4c7086c4",
   510 => x"c0c1029c",
   511 => x"eae4c287",
   512 => x"e149754a",
   513 => x"987087c9",
   514 => x"87f1c002",
   515 => x"49754a74",
   516 => x"efe14bcb",
   517 => x"02987087",
   518 => x"c087e2c0",
   519 => x"029c741e",
   520 => x"a6c487c7",
   521 => x"c578c048",
   522 => x"48a6c487",
   523 => x"66c478c1",
   524 => x"87eec949",
   525 => x"4c7086c4",
   526 => x"c0ff059c",
   527 => x"26487487",
   528 => x"0e87e7fc",
   529 => x"5d5c5b5e",
   530 => x"4b711e0e",
   531 => x"87c5059b",
   532 => x"e5c148c0",
   533 => x"4da3c887",
   534 => x"66d47dc0",
   535 => x"d487c702",
   536 => x"05bf9766",
   537 => x"48c087c5",
   538 => x"d487cfc1",
   539 => x"f3fd4966",
   540 => x"9c4c7087",
   541 => x"87c0c102",
   542 => x"6949a4dc",
   543 => x"49a4da7d",
   544 => x"9f4aa3c4",
   545 => x"e4c27a69",
   546 => x"d202bfe2",
   547 => x"49a4d487",
   548 => x"c049699f",
   549 => x"7199ffff",
   550 => x"7030d048",
   551 => x"c087c27e",
   552 => x"48496e7e",
   553 => x"7a70806a",
   554 => x"a3cc7bc0",
   555 => x"d0796a49",
   556 => x"79c049a3",
   557 => x"87c24874",
   558 => x"fa2648c0",
   559 => x"5e0e87ec",
   560 => x"0e5d5c5b",
   561 => x"f1c04c71",
   562 => x"78ff48f9",
   563 => x"c1029c74",
   564 => x"a4c887ca",
   565 => x"c1026949",
   566 => x"66d087c2",
   567 => x"82496c4a",
   568 => x"d05aa6d4",
   569 => x"c2b94d66",
   570 => x"4abfdee4",
   571 => x"9972baff",
   572 => x"c0029971",
   573 => x"a4c487e4",
   574 => x"f9496b4b",
   575 => x"7b7087f4",
   576 => x"bfdae4c2",
   577 => x"71816c49",
   578 => x"c2b9757c",
   579 => x"4abfdee4",
   580 => x"9972baff",
   581 => x"ff059971",
   582 => x"7c7587dc",
   583 => x"1e87cbf9",
   584 => x"4b711e73",
   585 => x"87c7029b",
   586 => x"6949a3c8",
   587 => x"c087c505",
   588 => x"87ebc048",
   589 => x"bff3e8c2",
   590 => x"49a3c44a",
   591 => x"89c24969",
   592 => x"bfdae4c2",
   593 => x"4aa27191",
   594 => x"bfdee4c2",
   595 => x"71996b49",
   596 => x"66c84aa2",
   597 => x"ea49721e",
   598 => x"86c487d2",
   599 => x"f8484970",
   600 => x"731e87cc",
   601 => x"9b4b711e",
   602 => x"c887c702",
   603 => x"056949a3",
   604 => x"48c087c5",
   605 => x"c287ebc0",
   606 => x"4abff3e8",
   607 => x"6949a3c4",
   608 => x"c289c249",
   609 => x"91bfdae4",
   610 => x"c24aa271",
   611 => x"49bfdee4",
   612 => x"a271996b",
   613 => x"1e66c84a",
   614 => x"c5e64972",
   615 => x"7086c487",
   616 => x"c9f74849",
   617 => x"5b5e0e87",
   618 => x"1e0e5d5c",
   619 => x"66d44b71",
   620 => x"732cc94c",
   621 => x"cfc1029b",
   622 => x"49a3c887",
   623 => x"c7c10269",
   624 => x"4da3d087",
   625 => x"c27d66d4",
   626 => x"49bfdee4",
   627 => x"4a6bb9ff",
   628 => x"ac717e99",
   629 => x"c087cd03",
   630 => x"a3cc7d7b",
   631 => x"49a3c44a",
   632 => x"87c2796a",
   633 => x"9c748c72",
   634 => x"4987dd02",
   635 => x"fb49731e",
   636 => x"86c487cc",
   637 => x"c74966d4",
   638 => x"cb0299ff",
   639 => x"dadcc287",
   640 => x"fc49731e",
   641 => x"86c487d9",
   642 => x"87def526",
   643 => x"711e731e",
   644 => x"c0029b4b",
   645 => x"e9c287e4",
   646 => x"4a735bc7",
   647 => x"e4c28ac2",
   648 => x"9249bfda",
   649 => x"bff3e8c2",
   650 => x"c2807248",
   651 => x"7158cbe9",
   652 => x"c230c448",
   653 => x"c058eae4",
   654 => x"e9c287ed",
   655 => x"e8c248c3",
   656 => x"c278bff7",
   657 => x"c248c7e9",
   658 => x"78bffbe8",
   659 => x"bfe2e4c2",
   660 => x"c287c902",
   661 => x"49bfdae4",
   662 => x"87c731c4",
   663 => x"bfffe8c2",
   664 => x"c231c449",
   665 => x"f459eae4",
   666 => x"5e0e87c4",
   667 => x"710e5c5b",
   668 => x"724bc04a",
   669 => x"e1c0029a",
   670 => x"49a2da87",
   671 => x"c24b699f",
   672 => x"02bfe2e4",
   673 => x"a2d487cf",
   674 => x"49699f49",
   675 => x"ffffc04c",
   676 => x"c234d09c",
   677 => x"744cc087",
   678 => x"4973b349",
   679 => x"f387edfd",
   680 => x"5e0e87ca",
   681 => x"0e5d5c5b",
   682 => x"4a7186f4",
   683 => x"9a727ec0",
   684 => x"c287d802",
   685 => x"c048d6dc",
   686 => x"cedcc278",
   687 => x"c7e9c248",
   688 => x"dcc278bf",
   689 => x"e9c248d2",
   690 => x"c278bfc3",
   691 => x"c048f7e4",
   692 => x"e6e4c250",
   693 => x"dcc249bf",
   694 => x"714abfd6",
   695 => x"ffc303aa",
   696 => x"cf497287",
   697 => x"e0c00599",
   698 => x"dadcc287",
   699 => x"cedcc21e",
   700 => x"dcc249bf",
   701 => x"a1c148ce",
   702 => x"efe37178",
   703 => x"c086c487",
   704 => x"c248f5f1",
   705 => x"cc78dadc",
   706 => x"f5f1c087",
   707 => x"e0c048bf",
   708 => x"f9f1c080",
   709 => x"d6dcc258",
   710 => x"80c148bf",
   711 => x"58dadcc2",
   712 => x"000c7527",
   713 => x"bf97bf00",
   714 => x"c2029d4d",
   715 => x"e5c387e2",
   716 => x"dbc202ad",
   717 => x"f5f1c087",
   718 => x"a3cb4bbf",
   719 => x"cf4c1149",
   720 => x"d2c105ac",
   721 => x"df497587",
   722 => x"cd89c199",
   723 => x"eae4c291",
   724 => x"4aa3c181",
   725 => x"a3c35112",
   726 => x"c551124a",
   727 => x"51124aa3",
   728 => x"124aa3c7",
   729 => x"4aa3c951",
   730 => x"a3ce5112",
   731 => x"d051124a",
   732 => x"51124aa3",
   733 => x"124aa3d2",
   734 => x"4aa3d451",
   735 => x"a3d65112",
   736 => x"d851124a",
   737 => x"51124aa3",
   738 => x"124aa3dc",
   739 => x"4aa3de51",
   740 => x"7ec15112",
   741 => x"7487f9c0",
   742 => x"0599c849",
   743 => x"7487eac0",
   744 => x"0599d049",
   745 => x"66dc87d0",
   746 => x"87cac002",
   747 => x"66dc4973",
   748 => x"0298700f",
   749 => x"056e87d3",
   750 => x"c287c6c0",
   751 => x"c048eae4",
   752 => x"f5f1c050",
   753 => x"e7c248bf",
   754 => x"f7e4c287",
   755 => x"7e50c048",
   756 => x"bfe6e4c2",
   757 => x"d6dcc249",
   758 => x"aa714abf",
   759 => x"87c1fc04",
   760 => x"bfc7e9c2",
   761 => x"87c8c005",
   762 => x"bfe2e4c2",
   763 => x"87fec102",
   764 => x"48f9f1c0",
   765 => x"dcc278ff",
   766 => x"ed49bfd2",
   767 => x"497087f4",
   768 => x"59d6dcc2",
   769 => x"c248a6c4",
   770 => x"78bfd2dc",
   771 => x"bfe2e4c2",
   772 => x"87d8c002",
   773 => x"cf4966c4",
   774 => x"f8ffffff",
   775 => x"c002a999",
   776 => x"4dc087c5",
   777 => x"c187e1c0",
   778 => x"87dcc04d",
   779 => x"cf4966c4",
   780 => x"a999f8ff",
   781 => x"87c8c002",
   782 => x"c048a6c8",
   783 => x"87c5c078",
   784 => x"c148a6c8",
   785 => x"4d66c878",
   786 => x"c0059d75",
   787 => x"66c487e0",
   788 => x"c289c249",
   789 => x"4abfdae4",
   790 => x"f3e8c291",
   791 => x"dcc24abf",
   792 => x"a17248ce",
   793 => x"d6dcc278",
   794 => x"f978c048",
   795 => x"48c087e3",
   796 => x"f5eb8ef4",
   797 => x"00000087",
   798 => x"ffffff00",
   799 => x"000c85ff",
   800 => x"000c8e00",
   801 => x"54414600",
   802 => x"20203233",
   803 => x"41460020",
   804 => x"20363154",
   805 => x"1e002020",
   806 => x"c348d4ff",
   807 => x"486878ff",
   808 => x"ff1e4f26",
   809 => x"ffc348d4",
   810 => x"48d0ff78",
   811 => x"ff78e1c8",
   812 => x"78d448d4",
   813 => x"48cbe9c2",
   814 => x"50bfd4ff",
   815 => x"ff1e4f26",
   816 => x"e0c048d0",
   817 => x"1e4f2678",
   818 => x"7087ccff",
   819 => x"c6029949",
   820 => x"a9fbc087",
   821 => x"7187f105",
   822 => x"0e4f2648",
   823 => x"0e5c5b5e",
   824 => x"4cc04b71",
   825 => x"7087f0fe",
   826 => x"c0029949",
   827 => x"ecc087f9",
   828 => x"f2c002a9",
   829 => x"a9fbc087",
   830 => x"87ebc002",
   831 => x"acb766cc",
   832 => x"d087c703",
   833 => x"87c20266",
   834 => x"99715371",
   835 => x"c187c202",
   836 => x"87c3fe84",
   837 => x"02994970",
   838 => x"ecc087cd",
   839 => x"87c702a9",
   840 => x"05a9fbc0",
   841 => x"d087d5ff",
   842 => x"87c30266",
   843 => x"c07b97c0",
   844 => x"c405a9ec",
   845 => x"c54a7487",
   846 => x"c04a7487",
   847 => x"48728a0a",
   848 => x"4d2687c2",
   849 => x"4b264c26",
   850 => x"fd1e4f26",
   851 => x"497087c9",
   852 => x"a9b7f0c0",
   853 => x"c087ca04",
   854 => x"01a9b7f9",
   855 => x"f0c087c3",
   856 => x"b7c1c189",
   857 => x"87ca04a9",
   858 => x"a9b7dac1",
   859 => x"c087c301",
   860 => x"487189f7",
   861 => x"5e0e4f26",
   862 => x"710e5c5b",
   863 => x"4cd4ff4a",
   864 => x"eac04972",
   865 => x"9b4b7087",
   866 => x"c187c202",
   867 => x"48d0ff8b",
   868 => x"c178c5c8",
   869 => x"49737cd5",
   870 => x"dac231c6",
   871 => x"4abf97de",
   872 => x"70b07148",
   873 => x"48d0ff7c",
   874 => x"487378c4",
   875 => x"0e87d5fe",
   876 => x"5d5c5b5e",
   877 => x"7186f80e",
   878 => x"fb7ec04c",
   879 => x"4bc087e4",
   880 => x"97dcf9c0",
   881 => x"a9c049bf",
   882 => x"fb87cf04",
   883 => x"83c187f9",
   884 => x"97dcf9c0",
   885 => x"06ab49bf",
   886 => x"f9c087f1",
   887 => x"02bf97dc",
   888 => x"f2fa87cf",
   889 => x"99497087",
   890 => x"c087c602",
   891 => x"f105a9ec",
   892 => x"fa4bc087",
   893 => x"4d7087e1",
   894 => x"c887dcfa",
   895 => x"d6fa58a6",
   896 => x"c14a7087",
   897 => x"49a4c883",
   898 => x"ad496997",
   899 => x"c087c702",
   900 => x"c005adff",
   901 => x"a4c987e7",
   902 => x"49699749",
   903 => x"02a966c4",
   904 => x"c04887c7",
   905 => x"d405a8ff",
   906 => x"49a4ca87",
   907 => x"aa496997",
   908 => x"c087c602",
   909 => x"c405aaff",
   910 => x"d07ec187",
   911 => x"adecc087",
   912 => x"c087c602",
   913 => x"c405adfb",
   914 => x"c14bc087",
   915 => x"fe026e7e",
   916 => x"e9f987e1",
   917 => x"f8487387",
   918 => x"87e6fb8e",
   919 => x"5b5e0e00",
   920 => x"1e0e5d5c",
   921 => x"4cc04b71",
   922 => x"c004ab4d",
   923 => x"f6c087e8",
   924 => x"9d751eef",
   925 => x"c087c402",
   926 => x"c187c24a",
   927 => x"f049724a",
   928 => x"86c487e0",
   929 => x"84c17e70",
   930 => x"87c2056e",
   931 => x"85c14c73",
   932 => x"ff06ac73",
   933 => x"486e87d8",
   934 => x"264d2626",
   935 => x"264b264c",
   936 => x"5b5e0e4f",
   937 => x"1e0e5d5c",
   938 => x"de494c71",
   939 => x"e5e9c291",
   940 => x"9785714d",
   941 => x"ddc1026d",
   942 => x"d0e9c287",
   943 => x"82744abf",
   944 => x"d8fe4972",
   945 => x"6e7e7087",
   946 => x"87f3c002",
   947 => x"4bd8e9c2",
   948 => x"49cb4a6e",
   949 => x"87d0c7ff",
   950 => x"93cb4b74",
   951 => x"83ceddc1",
   952 => x"fcc083c4",
   953 => x"49747bda",
   954 => x"87c9c3c1",
   955 => x"e9c27b75",
   956 => x"49bf97e4",
   957 => x"d8e9c21e",
   958 => x"e3ddc149",
   959 => x"7486c487",
   960 => x"f0c2c149",
   961 => x"c149c087",
   962 => x"c287cfc4",
   963 => x"c048cce9",
   964 => x"dd49c178",
   965 => x"fd2687cb",
   966 => x"6f4c87ff",
   967 => x"6e696461",
   968 => x"2e2e2e67",
   969 => x"5b5e0e00",
   970 => x"4b710e5c",
   971 => x"d0e9c24a",
   972 => x"497282bf",
   973 => x"7087e6fc",
   974 => x"c4029c4c",
   975 => x"e9ec4987",
   976 => x"d0e9c287",
   977 => x"c178c048",
   978 => x"87d5dc49",
   979 => x"0e87ccfd",
   980 => x"5d5c5b5e",
   981 => x"c286f40e",
   982 => x"c04ddadc",
   983 => x"48a6c44c",
   984 => x"e9c278c0",
   985 => x"c049bfd0",
   986 => x"c1c106a9",
   987 => x"dadcc287",
   988 => x"c0029848",
   989 => x"f6c087f8",
   990 => x"66c81eef",
   991 => x"c487c702",
   992 => x"78c048a6",
   993 => x"a6c487c5",
   994 => x"c478c148",
   995 => x"d1ec4966",
   996 => x"7086c487",
   997 => x"c484c14d",
   998 => x"80c14866",
   999 => x"c258a6c8",
  1000 => x"49bfd0e9",
  1001 => x"87c603ac",
  1002 => x"ff059d75",
  1003 => x"4cc087c8",
  1004 => x"c3029d75",
  1005 => x"f6c087e0",
  1006 => x"66c81eef",
  1007 => x"cc87c702",
  1008 => x"78c048a6",
  1009 => x"a6cc87c5",
  1010 => x"cc78c148",
  1011 => x"d1eb4966",
  1012 => x"7086c487",
  1013 => x"c2026e7e",
  1014 => x"496e87e9",
  1015 => x"699781cb",
  1016 => x"0299d049",
  1017 => x"c087d6c1",
  1018 => x"744ae5fc",
  1019 => x"c191cb49",
  1020 => x"7281cedd",
  1021 => x"c381c879",
  1022 => x"497451ff",
  1023 => x"e9c291de",
  1024 => x"85714de5",
  1025 => x"7d97c1c2",
  1026 => x"c049a5c1",
  1027 => x"e4c251e0",
  1028 => x"02bf97ea",
  1029 => x"84c187d2",
  1030 => x"c24ba5c2",
  1031 => x"db4aeae4",
  1032 => x"c3c2ff49",
  1033 => x"87dbc187",
  1034 => x"c049a5cd",
  1035 => x"c284c151",
  1036 => x"4a6e4ba5",
  1037 => x"c1ff49cb",
  1038 => x"c6c187ee",
  1039 => x"e1fac087",
  1040 => x"cb49744a",
  1041 => x"ceddc191",
  1042 => x"c2797281",
  1043 => x"bf97eae4",
  1044 => x"7487d802",
  1045 => x"c191de49",
  1046 => x"e5e9c284",
  1047 => x"c283714b",
  1048 => x"dd4aeae4",
  1049 => x"ffc0ff49",
  1050 => x"7487d887",
  1051 => x"c293de4b",
  1052 => x"cb83e5e9",
  1053 => x"51c049a3",
  1054 => x"6e7384c1",
  1055 => x"ff49cb4a",
  1056 => x"c487e5c0",
  1057 => x"80c14866",
  1058 => x"c758a6c8",
  1059 => x"c5c003ac",
  1060 => x"fc056e87",
  1061 => x"487487e0",
  1062 => x"fcf78ef4",
  1063 => x"1e731e87",
  1064 => x"cb494b71",
  1065 => x"ceddc191",
  1066 => x"4aa1c881",
  1067 => x"48dedac2",
  1068 => x"a1c95012",
  1069 => x"dcf9c04a",
  1070 => x"ca501248",
  1071 => x"e4e9c281",
  1072 => x"c2501148",
  1073 => x"bf97e4e9",
  1074 => x"49c01e49",
  1075 => x"87d0d6c1",
  1076 => x"48cce9c2",
  1077 => x"49c178de",
  1078 => x"2687c6d6",
  1079 => x"1e87fef6",
  1080 => x"cb494a71",
  1081 => x"ceddc191",
  1082 => x"1181c881",
  1083 => x"d0e9c248",
  1084 => x"d0e9c258",
  1085 => x"c178c048",
  1086 => x"87e5d549",
  1087 => x"c01e4f26",
  1088 => x"d5fcc049",
  1089 => x"1e4f2687",
  1090 => x"d2029971",
  1091 => x"e3dec187",
  1092 => x"f750c048",
  1093 => x"dfc3c180",
  1094 => x"c7ddc140",
  1095 => x"c187ce78",
  1096 => x"c148dfde",
  1097 => x"fc78c0dd",
  1098 => x"fec3c180",
  1099 => x"0e4f2678",
  1100 => x"0e5c5b5e",
  1101 => x"cb4a4c71",
  1102 => x"ceddc192",
  1103 => x"49a2c882",
  1104 => x"974ba2c9",
  1105 => x"971e4b6b",
  1106 => x"ca1e4969",
  1107 => x"c0491282",
  1108 => x"c087d0e7",
  1109 => x"87c9d449",
  1110 => x"f9c04974",
  1111 => x"8ef887d7",
  1112 => x"1e87f8f4",
  1113 => x"4b711e73",
  1114 => x"87c3ff49",
  1115 => x"fefe4973",
  1116 => x"87e9f487",
  1117 => x"711e731e",
  1118 => x"4aa3c64b",
  1119 => x"c187db02",
  1120 => x"87d6028a",
  1121 => x"dac1028a",
  1122 => x"c0028a87",
  1123 => x"028a87fc",
  1124 => x"8a87e1c0",
  1125 => x"c187cb02",
  1126 => x"49c787db",
  1127 => x"c187c0fd",
  1128 => x"e9c287de",
  1129 => x"c102bfd0",
  1130 => x"c14887cb",
  1131 => x"d4e9c288",
  1132 => x"87c1c158",
  1133 => x"bfd4e9c2",
  1134 => x"87f9c002",
  1135 => x"bfd0e9c2",
  1136 => x"c280c148",
  1137 => x"c058d4e9",
  1138 => x"e9c287eb",
  1139 => x"c649bfd0",
  1140 => x"d4e9c289",
  1141 => x"a9b7c059",
  1142 => x"c287da03",
  1143 => x"c048d0e9",
  1144 => x"c287d278",
  1145 => x"02bfd4e9",
  1146 => x"e9c287cb",
  1147 => x"c648bfd0",
  1148 => x"d4e9c280",
  1149 => x"d149c058",
  1150 => x"497387e7",
  1151 => x"87f5f6c0",
  1152 => x"0e87daf2",
  1153 => x"0e5c5b5e",
  1154 => x"66cc4c71",
  1155 => x"cb4b741e",
  1156 => x"ceddc193",
  1157 => x"4aa3c483",
  1158 => x"fafe496a",
  1159 => x"c2c187da",
  1160 => x"a3c87bdd",
  1161 => x"5166d449",
  1162 => x"d849a3c9",
  1163 => x"a3ca5166",
  1164 => x"5166dc49",
  1165 => x"87e3f126",
  1166 => x"5c5b5e0e",
  1167 => x"d0ff0e5d",
  1168 => x"59a6d886",
  1169 => x"c048a6c4",
  1170 => x"c180c478",
  1171 => x"c47866c4",
  1172 => x"c478c180",
  1173 => x"c278c180",
  1174 => x"c148d4e9",
  1175 => x"cce9c278",
  1176 => x"a8de48bf",
  1177 => x"f387cb05",
  1178 => x"497087e5",
  1179 => x"ce59a6c8",
  1180 => x"ede887f8",
  1181 => x"87cfe987",
  1182 => x"7087dce8",
  1183 => x"acfbc04c",
  1184 => x"87d0c102",
  1185 => x"c10566d4",
  1186 => x"1ec087c2",
  1187 => x"c11ec11e",
  1188 => x"c01ec1df",
  1189 => x"87ebfd49",
  1190 => x"4a66d0c1",
  1191 => x"496a82c4",
  1192 => x"517481c7",
  1193 => x"1ed81ec1",
  1194 => x"81c8496a",
  1195 => x"d887ece8",
  1196 => x"66c4c186",
  1197 => x"01a8c048",
  1198 => x"a6c487c7",
  1199 => x"ce78c148",
  1200 => x"66c4c187",
  1201 => x"cc88c148",
  1202 => x"87c358a6",
  1203 => x"cc87f8e7",
  1204 => x"78c248a6",
  1205 => x"cd029c74",
  1206 => x"66c487cc",
  1207 => x"66c8c148",
  1208 => x"c1cd03a8",
  1209 => x"48a6d887",
  1210 => x"eae678c0",
  1211 => x"c14c7087",
  1212 => x"c205acd0",
  1213 => x"66d887d6",
  1214 => x"87cee97e",
  1215 => x"a6dc4970",
  1216 => x"87d3e659",
  1217 => x"ecc04c70",
  1218 => x"eac105ac",
  1219 => x"4966c487",
  1220 => x"c0c191cb",
  1221 => x"a1c48166",
  1222 => x"c84d6a4a",
  1223 => x"66d84aa1",
  1224 => x"dfc3c152",
  1225 => x"87efe579",
  1226 => x"029c4c70",
  1227 => x"fbc087d8",
  1228 => x"87d202ac",
  1229 => x"dee55574",
  1230 => x"9c4c7087",
  1231 => x"c087c702",
  1232 => x"ff05acfb",
  1233 => x"e0c087ee",
  1234 => x"55c1c255",
  1235 => x"d47d97c0",
  1236 => x"a96e4966",
  1237 => x"c487db05",
  1238 => x"66c84866",
  1239 => x"87ca04a8",
  1240 => x"c14866c4",
  1241 => x"58a6c880",
  1242 => x"66c887c8",
  1243 => x"cc88c148",
  1244 => x"e2e458a6",
  1245 => x"c14c7087",
  1246 => x"c805acd0",
  1247 => x"4866d087",
  1248 => x"a6d480c1",
  1249 => x"acd0c158",
  1250 => x"87eafd02",
  1251 => x"d448a6dc",
  1252 => x"66d87866",
  1253 => x"a866dc48",
  1254 => x"87dcc905",
  1255 => x"48a6e0c0",
  1256 => x"c478f0c0",
  1257 => x"7866cc80",
  1258 => x"78c080c4",
  1259 => x"c048747e",
  1260 => x"f0c088fb",
  1261 => x"987058a6",
  1262 => x"87d7c802",
  1263 => x"c088cb48",
  1264 => x"7058a6f0",
  1265 => x"e9c00298",
  1266 => x"88c94887",
  1267 => x"58a6f0c0",
  1268 => x"c3029870",
  1269 => x"c44887e1",
  1270 => x"a6f0c088",
  1271 => x"02987058",
  1272 => x"c14887d6",
  1273 => x"a6f0c088",
  1274 => x"02987058",
  1275 => x"c787c8c3",
  1276 => x"e0c087db",
  1277 => x"78c048a6",
  1278 => x"c14866cc",
  1279 => x"58a6d080",
  1280 => x"7087d4e2",
  1281 => x"acecc04c",
  1282 => x"c087d502",
  1283 => x"c60266e0",
  1284 => x"a6e4c087",
  1285 => x"7487c95c",
  1286 => x"88f0c048",
  1287 => x"58a6e8c0",
  1288 => x"02acecc0",
  1289 => x"eee187cc",
  1290 => x"c04c7087",
  1291 => x"ff05acec",
  1292 => x"e0c087f4",
  1293 => x"66d41e66",
  1294 => x"ecc01e49",
  1295 => x"dfc11e66",
  1296 => x"66d41ec1",
  1297 => x"87fbf649",
  1298 => x"1eca1ec0",
  1299 => x"cb4966dc",
  1300 => x"66d8c191",
  1301 => x"48a6d881",
  1302 => x"d878a1c4",
  1303 => x"e149bf66",
  1304 => x"86d887f9",
  1305 => x"06a8b7c0",
  1306 => x"c187c7c1",
  1307 => x"c81ede1e",
  1308 => x"e149bf66",
  1309 => x"86c887e5",
  1310 => x"c0484970",
  1311 => x"e4c08808",
  1312 => x"b7c058a6",
  1313 => x"e9c006a8",
  1314 => x"66e0c087",
  1315 => x"a8b7dd48",
  1316 => x"6e87df03",
  1317 => x"e0c049bf",
  1318 => x"e0c08166",
  1319 => x"c1496651",
  1320 => x"81bf6e81",
  1321 => x"c051c1c2",
  1322 => x"c24966e0",
  1323 => x"81bf6e81",
  1324 => x"7ec151c0",
  1325 => x"e287dcc4",
  1326 => x"e4c087d0",
  1327 => x"c9e258a6",
  1328 => x"a6e8c087",
  1329 => x"a8ecc058",
  1330 => x"87cbc005",
  1331 => x"48a6e4c0",
  1332 => x"7866e0c0",
  1333 => x"ff87c4c0",
  1334 => x"c487fcde",
  1335 => x"91cb4966",
  1336 => x"4866c0c1",
  1337 => x"7e708071",
  1338 => x"82c84a6e",
  1339 => x"81ca496e",
  1340 => x"5166e0c0",
  1341 => x"4966e4c0",
  1342 => x"e0c081c1",
  1343 => x"48c18966",
  1344 => x"49703071",
  1345 => x"977189c1",
  1346 => x"c1edc27a",
  1347 => x"e0c049bf",
  1348 => x"6a972966",
  1349 => x"9871484a",
  1350 => x"58a6f0c0",
  1351 => x"81c4496e",
  1352 => x"66dc4d69",
  1353 => x"a866d848",
  1354 => x"87c8c002",
  1355 => x"c048a6d8",
  1356 => x"87c5c078",
  1357 => x"c148a6d8",
  1358 => x"1e66d878",
  1359 => x"751ee0c0",
  1360 => x"d6deff49",
  1361 => x"7086c887",
  1362 => x"acb7c04c",
  1363 => x"87d4c106",
  1364 => x"e0c08574",
  1365 => x"75897449",
  1366 => x"ded9c14b",
  1367 => x"edfe714a",
  1368 => x"85c287c6",
  1369 => x"4866e8c0",
  1370 => x"ecc080c1",
  1371 => x"ecc058a6",
  1372 => x"81c14966",
  1373 => x"c002a970",
  1374 => x"a6d887c8",
  1375 => x"c078c048",
  1376 => x"a6d887c5",
  1377 => x"d878c148",
  1378 => x"a4c21e66",
  1379 => x"48e0c049",
  1380 => x"49708871",
  1381 => x"ff49751e",
  1382 => x"c887c0dd",
  1383 => x"a8b7c086",
  1384 => x"87c0ff01",
  1385 => x"0266e8c0",
  1386 => x"6e87d1c0",
  1387 => x"c081c949",
  1388 => x"6e5166e8",
  1389 => x"efc4c148",
  1390 => x"87ccc078",
  1391 => x"81c9496e",
  1392 => x"486e51c2",
  1393 => x"78e3c5c1",
  1394 => x"c6c07ec1",
  1395 => x"f6dbff87",
  1396 => x"6e4c7087",
  1397 => x"87f5c002",
  1398 => x"c84866c4",
  1399 => x"c004a866",
  1400 => x"66c487cb",
  1401 => x"c880c148",
  1402 => x"e0c058a6",
  1403 => x"4866c887",
  1404 => x"a6cc88c1",
  1405 => x"87d5c058",
  1406 => x"05acc6c1",
  1407 => x"cc87c8c0",
  1408 => x"80c14866",
  1409 => x"ff58a6d0",
  1410 => x"7087fcda",
  1411 => x"4866d04c",
  1412 => x"a6d480c1",
  1413 => x"029c7458",
  1414 => x"c487cbc0",
  1415 => x"c8c14866",
  1416 => x"f204a866",
  1417 => x"daff87ff",
  1418 => x"66c487d4",
  1419 => x"03a8c748",
  1420 => x"c287e5c0",
  1421 => x"c048d4e9",
  1422 => x"4966c478",
  1423 => x"c0c191cb",
  1424 => x"a1c48166",
  1425 => x"c04a6a4a",
  1426 => x"66c47952",
  1427 => x"c880c148",
  1428 => x"a8c758a6",
  1429 => x"87dbff04",
  1430 => x"e08ed0ff",
  1431 => x"203a87fb",
  1432 => x"1e731e00",
  1433 => x"029b4b71",
  1434 => x"e9c287c6",
  1435 => x"78c048d0",
  1436 => x"e9c21ec7",
  1437 => x"1e49bfd0",
  1438 => x"1eceddc1",
  1439 => x"bfcce9c2",
  1440 => x"87f4ee49",
  1441 => x"e9c286cc",
  1442 => x"e949bfcc",
  1443 => x"9b7387f9",
  1444 => x"c187c802",
  1445 => x"c049cedd",
  1446 => x"ff87ece5",
  1447 => x"1e87fedf",
  1448 => x"48dedac2",
  1449 => x"dec150c0",
  1450 => x"c049bff1",
  1451 => x"c087c4fb",
  1452 => x"1e4f2648",
  1453 => x"c187e9c7",
  1454 => x"87e5fe49",
  1455 => x"87f1effe",
  1456 => x"cd029870",
  1457 => x"eef8fe87",
  1458 => x"02987087",
  1459 => x"4ac187c4",
  1460 => x"4ac087c2",
  1461 => x"ce059a72",
  1462 => x"c11ec087",
  1463 => x"c049c7dc",
  1464 => x"c487f3f0",
  1465 => x"c087fe86",
  1466 => x"c087ddff",
  1467 => x"d2dcc11e",
  1468 => x"e1f0c049",
  1469 => x"fe1ec087",
  1470 => x"497087e5",
  1471 => x"87d6f0c0",
  1472 => x"f887dcc3",
  1473 => x"534f268e",
  1474 => x"61662044",
  1475 => x"64656c69",
  1476 => x"6f42002e",
  1477 => x"6e69746f",
  1478 => x"2e2e2e67",
  1479 => x"e8c01e00",
  1480 => x"f3c087c1",
  1481 => x"87f687e6",
  1482 => x"c21e4f26",
  1483 => x"c048d0e9",
  1484 => x"cce9c278",
  1485 => x"fd78c048",
  1486 => x"87e187f9",
  1487 => x"4f2648c0",
  1488 => x"78452080",
  1489 => x"80007469",
  1490 => x"63614220",
  1491 => x"10df006b",
  1492 => x"2a650000",
  1493 => x"00000000",
  1494 => x"0010df00",
  1495 => x"002a8300",
  1496 => x"00000000",
  1497 => x"000010df",
  1498 => x"00002aa1",
  1499 => x"df000000",
  1500 => x"bf000010",
  1501 => x"0000002a",
  1502 => x"10df0000",
  1503 => x"2add0000",
  1504 => x"00000000",
  1505 => x"0010df00",
  1506 => x"002afb00",
  1507 => x"00000000",
  1508 => x"000010df",
  1509 => x"00002b19",
  1510 => x"df000000",
  1511 => x"00000010",
  1512 => x"00000000",
  1513 => x"11740000",
  1514 => x"00000000",
  1515 => x"00000000",
  1516 => x"0017b500",
  1517 => x"4f4f4200",
  1518 => x"20202054",
  1519 => x"4d4f5220",
  1520 => x"616f4c00",
  1521 => x"2e2a2064",
  1522 => x"f0fe1e00",
  1523 => x"cd78c048",
  1524 => x"26097909",
  1525 => x"fe1e1e4f",
  1526 => x"487ebff0",
  1527 => x"1e4f2626",
  1528 => x"c148f0fe",
  1529 => x"1e4f2678",
  1530 => x"c048f0fe",
  1531 => x"1e4f2678",
  1532 => x"52c04a71",
  1533 => x"0e4f2652",
  1534 => x"5d5c5b5e",
  1535 => x"7186f40e",
  1536 => x"7e6d974d",
  1537 => x"974ca5c1",
  1538 => x"a6c8486c",
  1539 => x"c4486e58",
  1540 => x"c505a866",
  1541 => x"c048ff87",
  1542 => x"caff87e6",
  1543 => x"49a5c287",
  1544 => x"714b6c97",
  1545 => x"6b974ba3",
  1546 => x"7e6c974b",
  1547 => x"80c1486e",
  1548 => x"c758a6c8",
  1549 => x"58a6cc98",
  1550 => x"fe7c9770",
  1551 => x"487387e1",
  1552 => x"4d268ef4",
  1553 => x"4b264c26",
  1554 => x"5e0e4f26",
  1555 => x"f40e5c5b",
  1556 => x"d84c7186",
  1557 => x"ffc34a66",
  1558 => x"4ba4c29a",
  1559 => x"73496c97",
  1560 => x"517249a1",
  1561 => x"6e7e6c97",
  1562 => x"c880c148",
  1563 => x"98c758a6",
  1564 => x"7058a6cc",
  1565 => x"ff8ef454",
  1566 => x"1e1e87ca",
  1567 => x"e087e8fd",
  1568 => x"c0494abf",
  1569 => x"0299c0e0",
  1570 => x"1e7287cb",
  1571 => x"49f7ecc2",
  1572 => x"c487f7fe",
  1573 => x"87fdfc86",
  1574 => x"c2fd7e70",
  1575 => x"4f262687",
  1576 => x"f7ecc21e",
  1577 => x"87c7fd49",
  1578 => x"49fae1c1",
  1579 => x"c587dafc",
  1580 => x"4f2687d9",
  1581 => x"5c5b5e0e",
  1582 => x"edc20e5d",
  1583 => x"c14abfd6",
  1584 => x"49bfc8e4",
  1585 => x"71bc724c",
  1586 => x"87dbfc4d",
  1587 => x"49744bc0",
  1588 => x"d50299d0",
  1589 => x"d0497587",
  1590 => x"c01e7199",
  1591 => x"daeac11e",
  1592 => x"1282734a",
  1593 => x"87e4c049",
  1594 => x"2cc186c8",
  1595 => x"abc8832d",
  1596 => x"87daff04",
  1597 => x"c187e8fb",
  1598 => x"c248c8e4",
  1599 => x"78bfd6ed",
  1600 => x"4c264d26",
  1601 => x"4f264b26",
  1602 => x"00000000",
  1603 => x"48d0ff1e",
  1604 => x"ff78e1c8",
  1605 => x"78c548d4",
  1606 => x"c30266c4",
  1607 => x"78e0c387",
  1608 => x"c60266c8",
  1609 => x"48d4ff87",
  1610 => x"ff78f0c3",
  1611 => x"787148d4",
  1612 => x"c848d0ff",
  1613 => x"e0c078e1",
  1614 => x"0e4f2678",
  1615 => x"0e5c5b5e",
  1616 => x"ecc24c71",
  1617 => x"eefa49f7",
  1618 => x"c04a7087",
  1619 => x"c204aab7",
  1620 => x"e0c387e3",
  1621 => x"87c905aa",
  1622 => x"48fee7c1",
  1623 => x"d4c278c1",
  1624 => x"aaf0c387",
  1625 => x"c187c905",
  1626 => x"c148fae7",
  1627 => x"87f5c178",
  1628 => x"bffee7c1",
  1629 => x"7287c702",
  1630 => x"b3c0c24b",
  1631 => x"4b7287c2",
  1632 => x"d1059c74",
  1633 => x"fae7c187",
  1634 => x"e7c11ebf",
  1635 => x"721ebffe",
  1636 => x"87f8fd49",
  1637 => x"e7c186c8",
  1638 => x"c002bffa",
  1639 => x"497387e0",
  1640 => x"9129b7c4",
  1641 => x"81dae9c1",
  1642 => x"9acf4a73",
  1643 => x"48c192c2",
  1644 => x"4a703072",
  1645 => x"4872baff",
  1646 => x"79709869",
  1647 => x"497387db",
  1648 => x"9129b7c4",
  1649 => x"81dae9c1",
  1650 => x"9acf4a73",
  1651 => x"48c392c2",
  1652 => x"4a703072",
  1653 => x"70b06948",
  1654 => x"fee7c179",
  1655 => x"c178c048",
  1656 => x"c048fae7",
  1657 => x"f7ecc278",
  1658 => x"87cbf849",
  1659 => x"b7c04a70",
  1660 => x"ddfd03aa",
  1661 => x"fc48c087",
  1662 => x"000087c8",
  1663 => x"00000000",
  1664 => x"711e0000",
  1665 => x"f2fc494a",
  1666 => x"1e4f2687",
  1667 => x"49724ac0",
  1668 => x"e9c191c4",
  1669 => x"79c081da",
  1670 => x"b7d082c1",
  1671 => x"87ee04aa",
  1672 => x"5e0e4f26",
  1673 => x"0e5d5c5b",
  1674 => x"faf64d71",
  1675 => x"c44a7587",
  1676 => x"c1922ab7",
  1677 => x"7582dae9",
  1678 => x"c29ccf4c",
  1679 => x"4b496a94",
  1680 => x"9bc32b74",
  1681 => x"307448c2",
  1682 => x"bcff4c70",
  1683 => x"98714874",
  1684 => x"caf67a70",
  1685 => x"fa487387",
  1686 => x"000087e6",
  1687 => x"80800000",
  1688 => x"80808080",
  1689 => x"80808080",
  1690 => x"80808080",
  1691 => x"80808080",
  1692 => x"80808080",
  1693 => x"80808080",
  1694 => x"80808080",
  1695 => x"80808080",
  1696 => x"80808080",
  1697 => x"80808080",
  1698 => x"80808080",
  1699 => x"80808080",
  1700 => x"80808080",
  1701 => x"80808080",
  1702 => x"1e168080",
  1703 => x"362e2526",
  1704 => x"ff1e3e3d",
  1705 => x"e1c848d0",
  1706 => x"ff487178",
  1707 => x"267808d4",
  1708 => x"d0ff1e4f",
  1709 => x"78e1c848",
  1710 => x"d4ff4871",
  1711 => x"66c47808",
  1712 => x"08d4ff48",
  1713 => x"1e4f2678",
  1714 => x"66c44a71",
  1715 => x"49721e49",
  1716 => x"ff87deff",
  1717 => x"e0c048d0",
  1718 => x"4f262678",
  1719 => x"c24a711e",
  1720 => x"c303aab7",
  1721 => x"87c28287",
  1722 => x"66c482ce",
  1723 => x"ff49721e",
  1724 => x"262687d5",
  1725 => x"d4ff1e4f",
  1726 => x"7affc34a",
  1727 => x"c848d0ff",
  1728 => x"7ade78e1",
  1729 => x"bfc1edc2",
  1730 => x"c848497a",
  1731 => x"717a7028",
  1732 => x"7028d048",
  1733 => x"d848717a",
  1734 => x"ff7a7028",
  1735 => x"e0c048d0",
  1736 => x"0e4f2678",
  1737 => x"5d5c5b5e",
  1738 => x"c24c710e",
  1739 => x"4dbfc1ed",
  1740 => x"d02b744b",
  1741 => x"83c19b66",
  1742 => x"04ab66d4",
  1743 => x"4bc087c2",
  1744 => x"66d04a74",
  1745 => x"ff317249",
  1746 => x"739975b9",
  1747 => x"70307248",
  1748 => x"b071484a",
  1749 => x"58c5edc2",
  1750 => x"2687dafe",
  1751 => x"264c264d",
  1752 => x"1e4f264b",
  1753 => x"c848d0ff",
  1754 => x"487178c9",
  1755 => x"7808d4ff",
  1756 => x"711e4f26",
  1757 => x"87eb494a",
  1758 => x"c848d0ff",
  1759 => x"1e4f2678",
  1760 => x"4b711e73",
  1761 => x"bfd1edc2",
  1762 => x"c287c302",
  1763 => x"d0ff87eb",
  1764 => x"78c9c848",
  1765 => x"e0c04973",
  1766 => x"48d4ffb1",
  1767 => x"edc27871",
  1768 => x"78c048c5",
  1769 => x"c50266c8",
  1770 => x"49ffc387",
  1771 => x"49c087c2",
  1772 => x"59cdedc2",
  1773 => x"c60266cc",
  1774 => x"d5d5c587",
  1775 => x"cf87c44a",
  1776 => x"c24affff",
  1777 => x"c25ad1ed",
  1778 => x"c148d1ed",
  1779 => x"2687c478",
  1780 => x"264c264d",
  1781 => x"0e4f264b",
  1782 => x"5d5c5b5e",
  1783 => x"c24a710e",
  1784 => x"4cbfcded",
  1785 => x"cb029a72",
  1786 => x"91c84987",
  1787 => x"4bf5edc1",
  1788 => x"87c48371",
  1789 => x"4bf5f1c1",
  1790 => x"49134dc0",
  1791 => x"edc29974",
  1792 => x"ffb9bfc9",
  1793 => x"787148d4",
  1794 => x"852cb7c1",
  1795 => x"04adb7c8",
  1796 => x"edc287e8",
  1797 => x"c848bfc5",
  1798 => x"c9edc280",
  1799 => x"87effe58",
  1800 => x"711e731e",
  1801 => x"9a4a134b",
  1802 => x"7287cb02",
  1803 => x"87e7fe49",
  1804 => x"059a4a13",
  1805 => x"dafe87f5",
  1806 => x"edc21e87",
  1807 => x"c249bfc5",
  1808 => x"c148c5ed",
  1809 => x"c0c478a1",
  1810 => x"db03a9b7",
  1811 => x"48d4ff87",
  1812 => x"bfc9edc2",
  1813 => x"c5edc278",
  1814 => x"edc249bf",
  1815 => x"a1c148c5",
  1816 => x"b7c0c478",
  1817 => x"87e504a9",
  1818 => x"c848d0ff",
  1819 => x"d1edc278",
  1820 => x"2678c048",
  1821 => x"0000004f",
  1822 => x"00000000",
  1823 => x"00000000",
  1824 => x"00005f5f",
  1825 => x"03030000",
  1826 => x"00030300",
  1827 => x"7f7f1400",
  1828 => x"147f7f14",
  1829 => x"2e240000",
  1830 => x"123a6b6b",
  1831 => x"366a4c00",
  1832 => x"32566c18",
  1833 => x"4f7e3000",
  1834 => x"683a7759",
  1835 => x"04000040",
  1836 => x"00000307",
  1837 => x"1c000000",
  1838 => x"0041633e",
  1839 => x"41000000",
  1840 => x"001c3e63",
  1841 => x"3e2a0800",
  1842 => x"2a3e1c1c",
  1843 => x"08080008",
  1844 => x"08083e3e",
  1845 => x"80000000",
  1846 => x"000060e0",
  1847 => x"08080000",
  1848 => x"08080808",
  1849 => x"00000000",
  1850 => x"00006060",
  1851 => x"30604000",
  1852 => x"03060c18",
  1853 => x"7f3e0001",
  1854 => x"3e7f4d59",
  1855 => x"06040000",
  1856 => x"00007f7f",
  1857 => x"63420000",
  1858 => x"464f5971",
  1859 => x"63220000",
  1860 => x"367f4949",
  1861 => x"161c1800",
  1862 => x"107f7f13",
  1863 => x"67270000",
  1864 => x"397d4545",
  1865 => x"7e3c0000",
  1866 => x"3079494b",
  1867 => x"01010000",
  1868 => x"070f7971",
  1869 => x"7f360000",
  1870 => x"367f4949",
  1871 => x"4f060000",
  1872 => x"1e3f6949",
  1873 => x"00000000",
  1874 => x"00006666",
  1875 => x"80000000",
  1876 => x"000066e6",
  1877 => x"08080000",
  1878 => x"22221414",
  1879 => x"14140000",
  1880 => x"14141414",
  1881 => x"22220000",
  1882 => x"08081414",
  1883 => x"03020000",
  1884 => x"060f5951",
  1885 => x"417f3e00",
  1886 => x"1e1f555d",
  1887 => x"7f7e0000",
  1888 => x"7e7f0909",
  1889 => x"7f7f0000",
  1890 => x"367f4949",
  1891 => x"3e1c0000",
  1892 => x"41414163",
  1893 => x"7f7f0000",
  1894 => x"1c3e6341",
  1895 => x"7f7f0000",
  1896 => x"41414949",
  1897 => x"7f7f0000",
  1898 => x"01010909",
  1899 => x"7f3e0000",
  1900 => x"7a7b4941",
  1901 => x"7f7f0000",
  1902 => x"7f7f0808",
  1903 => x"41000000",
  1904 => x"00417f7f",
  1905 => x"60200000",
  1906 => x"3f7f4040",
  1907 => x"087f7f00",
  1908 => x"4163361c",
  1909 => x"7f7f0000",
  1910 => x"40404040",
  1911 => x"067f7f00",
  1912 => x"7f7f060c",
  1913 => x"067f7f00",
  1914 => x"7f7f180c",
  1915 => x"7f3e0000",
  1916 => x"3e7f4141",
  1917 => x"7f7f0000",
  1918 => x"060f0909",
  1919 => x"417f3e00",
  1920 => x"407e7f61",
  1921 => x"7f7f0000",
  1922 => x"667f1909",
  1923 => x"6f260000",
  1924 => x"327b594d",
  1925 => x"01010000",
  1926 => x"01017f7f",
  1927 => x"7f3f0000",
  1928 => x"3f7f4040",
  1929 => x"3f0f0000",
  1930 => x"0f3f7070",
  1931 => x"307f7f00",
  1932 => x"7f7f3018",
  1933 => x"36634100",
  1934 => x"63361c1c",
  1935 => x"06030141",
  1936 => x"03067c7c",
  1937 => x"59716101",
  1938 => x"4143474d",
  1939 => x"7f000000",
  1940 => x"0041417f",
  1941 => x"06030100",
  1942 => x"6030180c",
  1943 => x"41000040",
  1944 => x"007f7f41",
  1945 => x"060c0800",
  1946 => x"080c0603",
  1947 => x"80808000",
  1948 => x"80808080",
  1949 => x"00000000",
  1950 => x"00040703",
  1951 => x"74200000",
  1952 => x"787c5454",
  1953 => x"7f7f0000",
  1954 => x"387c4444",
  1955 => x"7c380000",
  1956 => x"00444444",
  1957 => x"7c380000",
  1958 => x"7f7f4444",
  1959 => x"7c380000",
  1960 => x"185c5454",
  1961 => x"7e040000",
  1962 => x"0005057f",
  1963 => x"bc180000",
  1964 => x"7cfca4a4",
  1965 => x"7f7f0000",
  1966 => x"787c0404",
  1967 => x"00000000",
  1968 => x"00407d3d",
  1969 => x"80800000",
  1970 => x"007dfd80",
  1971 => x"7f7f0000",
  1972 => x"446c3810",
  1973 => x"00000000",
  1974 => x"00407f3f",
  1975 => x"0c7c7c00",
  1976 => x"787c0c18",
  1977 => x"7c7c0000",
  1978 => x"787c0404",
  1979 => x"7c380000",
  1980 => x"387c4444",
  1981 => x"fcfc0000",
  1982 => x"183c2424",
  1983 => x"3c180000",
  1984 => x"fcfc2424",
  1985 => x"7c7c0000",
  1986 => x"080c0404",
  1987 => x"5c480000",
  1988 => x"20745454",
  1989 => x"3f040000",
  1990 => x"0044447f",
  1991 => x"7c3c0000",
  1992 => x"7c7c4040",
  1993 => x"3c1c0000",
  1994 => x"1c3c6060",
  1995 => x"607c3c00",
  1996 => x"3c7c6030",
  1997 => x"386c4400",
  1998 => x"446c3810",
  1999 => x"bc1c0000",
  2000 => x"1c3c60e0",
  2001 => x"64440000",
  2002 => x"444c5c74",
  2003 => x"08080000",
  2004 => x"4141773e",
  2005 => x"00000000",
  2006 => x"00007f7f",
  2007 => x"41410000",
  2008 => x"08083e77",
  2009 => x"01010200",
  2010 => x"01020203",
  2011 => x"7f7f7f00",
  2012 => x"7f7f7f7f",
  2013 => x"1c080800",
  2014 => x"7f3e3e1c",
  2015 => x"3e7f7f7f",
  2016 => x"081c1c3e",
  2017 => x"18100008",
  2018 => x"10187c7c",
  2019 => x"30100000",
  2020 => x"10307c7c",
  2021 => x"60301000",
  2022 => x"061e7860",
  2023 => x"3c664200",
  2024 => x"42663c18",
  2025 => x"6a387800",
  2026 => x"386cc6c2",
  2027 => x"00006000",
  2028 => x"60000060",
  2029 => x"5b5e0e00",
  2030 => x"1e0e5d5c",
  2031 => x"edc24c71",
  2032 => x"c04dbfe2",
  2033 => x"741ec04b",
  2034 => x"87c702ab",
  2035 => x"c048a6c4",
  2036 => x"c487c578",
  2037 => x"78c148a6",
  2038 => x"731e66c4",
  2039 => x"87dfee49",
  2040 => x"e0c086c8",
  2041 => x"87efef49",
  2042 => x"6a4aa5c4",
  2043 => x"87f0f049",
  2044 => x"cb87c6f1",
  2045 => x"c883c185",
  2046 => x"ff04abb7",
  2047 => x"262687c7",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
