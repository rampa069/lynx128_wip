library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom2 is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"264c264d",
     1 => x"1e4f264b",
     2 => x"edc24a71",
     3 => x"edc25ae6",
     4 => x"78c748e6",
     5 => x"87ddfe49",
     6 => x"731e4f26",
     7 => x"c04a711e",
     8 => x"d303aab7",
     9 => x"ebcdc287",
    10 => x"87c405bf",
    11 => x"87c24bc1",
    12 => x"cdc24bc0",
    13 => x"87c45bef",
    14 => x"5aefcdc2",
    15 => x"bfebcdc2",
    16 => x"c19ac14a",
    17 => x"ec49a2c0",
    18 => x"48fc87e8",
    19 => x"bfebcdc2",
    20 => x"87effe78",
    21 => x"c44a711e",
    22 => x"49721e66",
    23 => x"2687fde9",
    24 => x"c21e4f26",
    25 => x"49bfebcd",
    26 => x"c287d7e6",
    27 => x"e848daed",
    28 => x"edc278bf",
    29 => x"bfec48d6",
    30 => x"daedc278",
    31 => x"c3494abf",
    32 => x"b7c899ff",
    33 => x"7148722a",
    34 => x"e2edc2b0",
    35 => x"0e4f2658",
    36 => x"5d5c5b5e",
    37 => x"ff4b710e",
    38 => x"edc287c8",
    39 => x"50c048d5",
    40 => x"fde54973",
    41 => x"4c497087",
    42 => x"eecb9cc2",
    43 => x"87c3cb49",
    44 => x"c24d4970",
    45 => x"bf97d5ed",
    46 => x"87e2c105",
    47 => x"c24966d0",
    48 => x"99bfdeed",
    49 => x"d487d605",
    50 => x"edc24966",
    51 => x"0599bfd6",
    52 => x"497387cb",
    53 => x"7087cbe5",
    54 => x"c1c10298",
    55 => x"fe4cc187",
    56 => x"497587c0",
    57 => x"7087d8ca",
    58 => x"87c60298",
    59 => x"48d5edc2",
    60 => x"edc250c1",
    61 => x"05bf97d5",
    62 => x"c287e3c0",
    63 => x"49bfdeed",
    64 => x"059966d0",
    65 => x"c287d6ff",
    66 => x"49bfd6ed",
    67 => x"059966d4",
    68 => x"7387caff",
    69 => x"87cae449",
    70 => x"fe059870",
    71 => x"487487ff",
    72 => x"0e87dcfb",
    73 => x"5d5c5b5e",
    74 => x"c086f40e",
    75 => x"bfec4c4d",
    76 => x"48a6c47e",
    77 => x"bfe2edc2",
    78 => x"c01ec178",
    79 => x"fd49c71e",
    80 => x"86c887cd",
    81 => x"cd029870",
    82 => x"fb49ff87",
    83 => x"dac187cc",
    84 => x"87cee349",
    85 => x"edc24dc1",
    86 => x"02bf97d5",
    87 => x"fed487c3",
    88 => x"daedc287",
    89 => x"cdc24bbf",
    90 => x"c005bfeb",
    91 => x"fdc387e9",
    92 => x"87eee249",
    93 => x"e249fac3",
    94 => x"497387e8",
    95 => x"7199ffc3",
    96 => x"fb49c01e",
    97 => x"497387ce",
    98 => x"7129b7c8",
    99 => x"fb49c11e",
   100 => x"86c887c2",
   101 => x"c287fac5",
   102 => x"4bbfdeed",
   103 => x"87dd029b",
   104 => x"bfe7cdc2",
   105 => x"87d7c749",
   106 => x"c4059870",
   107 => x"d24bc087",
   108 => x"49e0c287",
   109 => x"c287fcc6",
   110 => x"c658ebcd",
   111 => x"e7cdc287",
   112 => x"7378c048",
   113 => x"0599c249",
   114 => x"ebc387cd",
   115 => x"87d2e149",
   116 => x"99c24970",
   117 => x"fb87c202",
   118 => x"c149734c",
   119 => x"87cd0599",
   120 => x"e049f4c3",
   121 => x"497087fc",
   122 => x"c20299c2",
   123 => x"734cfa87",
   124 => x"0599c849",
   125 => x"f5c387cd",
   126 => x"87e6e049",
   127 => x"99c24970",
   128 => x"c287d402",
   129 => x"02bfe6ed",
   130 => x"c14887c9",
   131 => x"eaedc288",
   132 => x"ff87c258",
   133 => x"734dc14c",
   134 => x"0599c449",
   135 => x"f2c387ce",
   136 => x"fddfff49",
   137 => x"c2497087",
   138 => x"87db0299",
   139 => x"bfe6edc2",
   140 => x"b7c7487e",
   141 => x"87cb03a8",
   142 => x"80c1486e",
   143 => x"58eaedc2",
   144 => x"fe87c2c0",
   145 => x"c34dc14c",
   146 => x"dfff49fd",
   147 => x"497087d4",
   148 => x"d50299c2",
   149 => x"e6edc287",
   150 => x"c9c002bf",
   151 => x"e6edc287",
   152 => x"c078c048",
   153 => x"4cfd87c2",
   154 => x"fac34dc1",
   155 => x"f1deff49",
   156 => x"c2497087",
   157 => x"87d90299",
   158 => x"bfe6edc2",
   159 => x"a8b7c748",
   160 => x"87c9c003",
   161 => x"48e6edc2",
   162 => x"c2c078c7",
   163 => x"c14cfc87",
   164 => x"acb7c04d",
   165 => x"87d1c003",
   166 => x"c14a66c4",
   167 => x"026a82d8",
   168 => x"6a87c6c0",
   169 => x"7349744b",
   170 => x"c31ec00f",
   171 => x"dac11ef0",
   172 => x"87dbf749",
   173 => x"987086c8",
   174 => x"87e2c002",
   175 => x"c248a6c8",
   176 => x"78bfe6ed",
   177 => x"cb4966c8",
   178 => x"4866c491",
   179 => x"7e708071",
   180 => x"c002bf6e",
   181 => x"bf6e87c8",
   182 => x"4966c84b",
   183 => x"9d750f73",
   184 => x"87c8c002",
   185 => x"bfe6edc2",
   186 => x"87c9f349",
   187 => x"bfefcdc2",
   188 => x"87ddc002",
   189 => x"87c7c249",
   190 => x"c0029870",
   191 => x"edc287d3",
   192 => x"f249bfe6",
   193 => x"49c087ef",
   194 => x"c287cff4",
   195 => x"c048efcd",
   196 => x"f38ef478",
   197 => x"5e0e87e9",
   198 => x"0e5d5c5b",
   199 => x"c24c711e",
   200 => x"49bfe2ed",
   201 => x"4da1cdc1",
   202 => x"6981d1c1",
   203 => x"029c747e",
   204 => x"a5c487cf",
   205 => x"c27b744b",
   206 => x"49bfe2ed",
   207 => x"6e87c8f3",
   208 => x"059c747b",
   209 => x"4bc087c4",
   210 => x"4bc187c2",
   211 => x"c9f34973",
   212 => x"0266d487",
   213 => x"da4987c7",
   214 => x"c24a7087",
   215 => x"c24ac087",
   216 => x"265af3cd",
   217 => x"0087d8f2",
   218 => x"00000000",
   219 => x"00000000",
   220 => x"1e000000",
   221 => x"c8ff4a71",
   222 => x"a17249bf",
   223 => x"1e4f2648",
   224 => x"89bfc8ff",
   225 => x"c0c0c0c2",
   226 => x"01a9c0c0",
   227 => x"4ac087c4",
   228 => x"4ac187c2",
   229 => x"4f264872",
   230 => x"5c5b5e0e",
   231 => x"4b710e5d",
   232 => x"d04cd4ff",
   233 => x"78c04866",
   234 => x"dbff49d6",
   235 => x"ffc387f4",
   236 => x"c3496c7c",
   237 => x"4d7199ff",
   238 => x"99f0c349",
   239 => x"05a9e0c1",
   240 => x"ffc387cb",
   241 => x"c3486c7c",
   242 => x"0866d098",
   243 => x"7cffc378",
   244 => x"c8494a6c",
   245 => x"7cffc331",
   246 => x"b2714a6c",
   247 => x"31c84972",
   248 => x"6c7cffc3",
   249 => x"72b2714a",
   250 => x"c331c849",
   251 => x"4a6c7cff",
   252 => x"d0ffb271",
   253 => x"78e0c048",
   254 => x"c2029b73",
   255 => x"757b7287",
   256 => x"264d2648",
   257 => x"264b264c",
   258 => x"4f261e4f",
   259 => x"5c5b5e0e",
   260 => x"7686f80e",
   261 => x"49a6c81e",
   262 => x"c487fdfd",
   263 => x"6e4b7086",
   264 => x"01a8c048",
   265 => x"7387c6c3",
   266 => x"9af0c34a",
   267 => x"02aad0c1",
   268 => x"e0c187c7",
   269 => x"f4c205aa",
   270 => x"c8497387",
   271 => x"87c30299",
   272 => x"7387c6ff",
   273 => x"c29cc34c",
   274 => x"cdc105ac",
   275 => x"4966c487",
   276 => x"1e7131c9",
   277 => x"d44a66c4",
   278 => x"eaedc292",
   279 => x"fe817249",
   280 => x"c487c2d5",
   281 => x"c01e4966",
   282 => x"d9ff49e3",
   283 => x"49d887d9",
   284 => x"87eed8ff",
   285 => x"c21ec0c8",
   286 => x"fd49dadc",
   287 => x"ff87d7f1",
   288 => x"e0c048d0",
   289 => x"dadcc278",
   290 => x"4a66d01e",
   291 => x"edc292d4",
   292 => x"817249ea",
   293 => x"87cad3fe",
   294 => x"acc186d0",
   295 => x"87cdc105",
   296 => x"c94966c4",
   297 => x"c41e7131",
   298 => x"92d44a66",
   299 => x"49eaedc2",
   300 => x"d3fe8172",
   301 => x"dcc287ef",
   302 => x"66c81eda",
   303 => x"c292d44a",
   304 => x"7249eaed",
   305 => x"d6d1fe81",
   306 => x"4966c887",
   307 => x"49e3c01e",
   308 => x"87f3d7ff",
   309 => x"d7ff49d7",
   310 => x"c0c887c8",
   311 => x"dadcc21e",
   312 => x"e0effd49",
   313 => x"ff86d087",
   314 => x"e0c048d0",
   315 => x"fc8ef878",
   316 => x"5e0e87d1",
   317 => x"0e5d5c5b",
   318 => x"ff4d711e",
   319 => x"66d44cd4",
   320 => x"b7c3487e",
   321 => x"87c506a8",
   322 => x"e2c148c0",
   323 => x"fe497587",
   324 => x"7587e3e1",
   325 => x"4b66c41e",
   326 => x"edc293d4",
   327 => x"497383ea",
   328 => x"87dfccfe",
   329 => x"4b6b83c8",
   330 => x"c848d0ff",
   331 => x"7cdd78e1",
   332 => x"ffc34973",
   333 => x"737c7199",
   334 => x"29b7c849",
   335 => x"7199ffc3",
   336 => x"d049737c",
   337 => x"ffc329b7",
   338 => x"737c7199",
   339 => x"29b7d849",
   340 => x"7cc07c71",
   341 => x"7c7c7c7c",
   342 => x"7c7c7c7c",
   343 => x"c07c7c7c",
   344 => x"66c478e0",
   345 => x"ff49dc1e",
   346 => x"c887dcd5",
   347 => x"26487386",
   348 => x"0e87cefa",
   349 => x"5d5c5b5e",
   350 => x"7e711e0e",
   351 => x"6e4bd4ff",
   352 => x"feedc21e",
   353 => x"facafe49",
   354 => x"7086c487",
   355 => x"c3029d4d",
   356 => x"eec287c3",
   357 => x"6e4cbfc6",
   358 => x"d9dffe49",
   359 => x"48d0ff87",
   360 => x"c178c5c8",
   361 => x"4ac07bd6",
   362 => x"82c17b15",
   363 => x"aab7e0c0",
   364 => x"ff87f504",
   365 => x"78c448d0",
   366 => x"c178c5c8",
   367 => x"7bc17bd3",
   368 => x"9c7478c4",
   369 => x"87fcc102",
   370 => x"7edadcc2",
   371 => x"8c4dc0c8",
   372 => x"03acb7c0",
   373 => x"c0c887c6",
   374 => x"4cc04da4",
   375 => x"97cbe9c2",
   376 => x"99d049bf",
   377 => x"c087d202",
   378 => x"feedc21e",
   379 => x"eeccfe49",
   380 => x"7086c487",
   381 => x"efc04a49",
   382 => x"dadcc287",
   383 => x"feedc21e",
   384 => x"daccfe49",
   385 => x"7086c487",
   386 => x"d0ff4a49",
   387 => x"78c5c848",
   388 => x"6e7bd4c1",
   389 => x"6e7bbf97",
   390 => x"7080c148",
   391 => x"058dc17e",
   392 => x"ff87f0ff",
   393 => x"78c448d0",
   394 => x"c5059a72",
   395 => x"c048c087",
   396 => x"1ec187e5",
   397 => x"49feedc2",
   398 => x"87c2cafe",
   399 => x"9c7486c4",
   400 => x"87c4fe05",
   401 => x"c848d0ff",
   402 => x"d3c178c5",
   403 => x"c47bc07b",
   404 => x"c248c178",
   405 => x"2648c087",
   406 => x"4c264d26",
   407 => x"4f264b26",
   408 => x"5c5b5e0e",
   409 => x"cc4b710e",
   410 => x"87d80266",
   411 => x"8cf0c04c",
   412 => x"7487d802",
   413 => x"028ac14a",
   414 => x"028a87d1",
   415 => x"028a87cd",
   416 => x"87d787c9",
   417 => x"eafb4973",
   418 => x"7487d087",
   419 => x"f949c01e",
   420 => x"1e7487e0",
   421 => x"d9f94973",
   422 => x"fe86c887",
   423 => x"1e0087fc",
   424 => x"bfeddbc2",
   425 => x"c2b9c149",
   426 => x"ff59f1db",
   427 => x"ffc348d4",
   428 => x"48d0ff78",
   429 => x"ff78e1c8",
   430 => x"78c148d4",
   431 => x"787131c4",
   432 => x"c048d0ff",
   433 => x"4f2678e0",
   434 => x"e1dbc21e",
   435 => x"feedc21e",
   436 => x"eec5fe49",
   437 => x"7086c487",
   438 => x"87c30298",
   439 => x"2687c0ff",
   440 => x"4b35314f",
   441 => x"20205a48",
   442 => x"47464320",
   443 => x"00000000",
   444 => x"00000000",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
