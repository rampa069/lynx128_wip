//-------------------------------------------------------------------------------------------------
module digit2 #
//-------------------------------------------------------------------------------------------------
(
	parameter X = 0,
	parameter Y = 0
)
//-------------------------------------------------------------------------------------------------
(
	input  wire       clock,
	input  wire       ce,
	input  wire       hs,
	input  wire       vs,
	input  wire[ 7:0] value,
	output wire       pixel,
	output wire       de
);
//-------------------------------------------------------------------------------------------------

reg[7:0] font[127:0];
initial
begin
font['h00] = 8'b000000000; font['h08] = 8'b000000000; font['h10] = 8'b000000000; font['h18] = 8'b000000000;
font['h01] = 8'b001111100; font['h09] = 8'b000011000; font['h11] = 8'b001111100; font['h19] = 8'b011111100;
font['h02] = 8'b011000110; font['h0A] = 8'b000111000; font['h12] = 8'b000000110; font['h1A] = 8'b000000110;
font['h03] = 8'b011010110; font['h0B] = 8'b001111000; font['h13] = 8'b000000110; font['h1B] = 8'b000000110;
font['h04] = 8'b011010110; font['h0C] = 8'b000011000; font['h14] = 8'b001111100; font['h1C] = 8'b001111100;
font['h05] = 8'b011010110; font['h0D] = 8'b000011000; font['h15] = 8'b011000000; font['h1D] = 8'b000000110;
font['h06] = 8'b011000110; font['h0E] = 8'b000011000; font['h16] = 8'b011000000; font['h1E] = 8'b000000110;
font['h07] = 8'b001111100; font['h0F] = 8'b000011000; font['h17] = 8'b011111110; font['h1F] = 8'b011111100;

font['h20] = 8'b000000000; font['h28] = 8'b000000000; font['h30] = 8'b000000000; font['h38] = 8'b000000000;
font['h21] = 8'b011000000; font['h29] = 8'b011111100; font['h31] = 8'b001111100; font['h39] = 8'b011111110;
font['h22] = 8'b011000000; font['h2A] = 8'b011000000; font['h32] = 8'b011000000; font['h3A] = 8'b000000110;
font['h23] = 8'b011000000; font['h2B] = 8'b011000000; font['h33] = 8'b011000000; font['h3B] = 8'b000001100;
font['h24] = 8'b011001100; font['h2C] = 8'b011111100; font['h34] = 8'b011111100; font['h3C] = 8'b000011000;
font['h25] = 8'b011111110; font['h2D] = 8'b000000110; font['h35] = 8'b011000110; font['h3D] = 8'b000110000;
font['h26] = 8'b000001100; font['h2E] = 8'b000000110; font['h36] = 8'b011000110; font['h3E] = 8'b000110000;
font['h27] = 8'b000001100; font['h2F] = 8'b011111100; font['h37] = 8'b001111100; font['h3F] = 8'b000110000;

font['h40] = 8'b000000000; font['h48] = 8'b000000000; font['h50] = 8'b000000000; font['h58] = 8'b000000000;
font['h41] = 8'b001111100; font['h49] = 8'b001111100; font['h51] = 8'b001111100; font['h59] = 8'b011111100;
font['h42] = 8'b011000110; font['h4A] = 8'b011000110; font['h52] = 8'b011000110; font['h5A] = 8'b011000110;
font['h43] = 8'b011000110; font['h4B] = 8'b011000110; font['h53] = 8'b011000110; font['h5B] = 8'b011000110;
font['h44] = 8'b001111100; font['h4C] = 8'b001111110; font['h54] = 8'b011111110; font['h5C] = 8'b011111100;
font['h45] = 8'b011000110; font['h4D] = 8'b000000110; font['h55] = 8'b011000110; font['h5D] = 8'b011000110;
font['h46] = 8'b011000110; font['h4E] = 8'b000000110; font['h56] = 8'b011000110; font['h5E] = 8'b011000110;
font['h47] = 8'b001111100; font['h4F] = 8'b001111100; font['h57] = 8'b011000110; font['h5F] = 8'b011111100;

font['h60] = 8'b000000000; font['h68] = 8'b000000000; font['h70] = 8'b000000000; font['h78] = 8'b000000000;
font['h61] = 8'b001111110; font['h69] = 8'b011111100; font['h71] = 8'b011111110; font['h79] = 8'b011111110;
font['h62] = 8'b011000000; font['h6A] = 8'b011000110; font['h72] = 8'b011000000; font['h7A] = 8'b011000000;
font['h63] = 8'b011000000; font['h6B] = 8'b011000110; font['h73] = 8'b011000000; font['h7B] = 8'b011000000;
font['h64] = 8'b011000000; font['h6C] = 8'b011000110; font['h74] = 8'b011111100; font['h7C] = 8'b011111100;
font['h65] = 8'b011000000; font['h6D] = 8'b011000110; font['h75] = 8'b011000000; font['h7D] = 8'b011000000;
font['h66] = 8'b011000000; font['h6E] = 8'b011000110; font['h76] = 8'b011000000; font['h7E] = 8'b011000000;
font['h67] = 8'b001111110; font['h6F] = 8'b011111100; font['h77] = 8'b011111110; font['h7F] = 8'b011000000;
end

//-------------------------------------------------------------------------------------------------

reg vsd;
reg yrs;
always @(posedge clock) if(ce) begin vsd <= vs; yrs <= ~vs&vsd; end

reg hsd;
reg xrs;
always @(posedge clock) if(ce) begin hsd <= hs; xrs <= ~hs&hsd; end

reg[9:0] y;
always @(posedge clock) if(ce) if(yrs) y <= 1'd0; else if(xrs) y <= y+1'd1;

reg[9:0] x;
always @(posedge clock) if(ce) if(xrs) x <= 1'd0; else x <= x+1'd1;

reg iy;
reg ix;
reg[2:0] yc;
reg[3:0] xc;
reg[7:0] bmp;
always @(posedge clock) if(ce)
begin
	if(y == Y) iy <= 1'b1;
	if(x == X) if(iy) ix <= 1'b1;

	if(ix)
	begin
		xc <= xc+1'd1;
		if(xc[2:0] == 0) bmp <= font[{ xc[3] ? value[3:0] : value[7:4], yc }]; else bmp <= { bmp[6:0], 1'b0 };

		if(xc == 15)
		begin
			yc <= yc+1'd1;
			ix <= 1'b0;

			if(yc == 7) iy <= 1'b0;
		end
	end
end

assign pixel = bmp[7];
assign de = ix && iy;

//-------------------------------------------------------------------------------------------------
endmodule
//-------------------------------------------------------------------------------------------------
